library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"dcefc287",
    12 => x"86c0c64e",
    13 => x"49dcefc2",
    14 => x"48e8dcc2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087cbdc",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"48111e4f",
    50 => x"7808d4ff",
    51 => x"c14866c4",
    52 => x"58a6c888",
    53 => x"ed059870",
    54 => x"1e4f2687",
    55 => x"c348d4ff",
    56 => x"516878ff",
    57 => x"c14866c4",
    58 => x"58a6c888",
    59 => x"eb059870",
    60 => x"1e4f2687",
    61 => x"d4ff1e73",
    62 => x"7bffc34b",
    63 => x"ffc34a6b",
    64 => x"c8496b7b",
    65 => x"c3b17232",
    66 => x"4a6b7bff",
    67 => x"b27131c8",
    68 => x"6b7bffc3",
    69 => x"7232c849",
    70 => x"c44871b1",
    71 => x"264d2687",
    72 => x"264b264c",
    73 => x"5b5e0e4f",
    74 => x"710e5d5c",
    75 => x"4cd4ff4a",
    76 => x"ffc34972",
    77 => x"c27c7199",
    78 => x"05bfe8dc",
    79 => x"66d087c8",
    80 => x"d430c948",
    81 => x"66d058a6",
    82 => x"c329d849",
    83 => x"7c7199ff",
    84 => x"d04966d0",
    85 => x"99ffc329",
    86 => x"66d07c71",
    87 => x"c329c849",
    88 => x"7c7199ff",
    89 => x"c34966d0",
    90 => x"7c7199ff",
    91 => x"29d04972",
    92 => x"7199ffc3",
    93 => x"c94b6c7c",
    94 => x"c34dfff0",
    95 => x"d005abff",
    96 => x"7cffc387",
    97 => x"8dc14b6c",
    98 => x"c387c602",
    99 => x"f002abff",
   100 => x"fe487387",
   101 => x"c01e87c7",
   102 => x"48d4ff49",
   103 => x"c178ffc3",
   104 => x"b7c8c381",
   105 => x"87f104a9",
   106 => x"731e4f26",
   107 => x"c487e71e",
   108 => x"c04bdff8",
   109 => x"f0ffc01e",
   110 => x"fd49f7c1",
   111 => x"86c487e7",
   112 => x"c005a8c1",
   113 => x"d4ff87ea",
   114 => x"78ffc348",
   115 => x"c0c0c0c1",
   116 => x"c01ec0c0",
   117 => x"e9c1f0e1",
   118 => x"87c9fd49",
   119 => x"987086c4",
   120 => x"ff87ca05",
   121 => x"ffc348d4",
   122 => x"cb48c178",
   123 => x"87e6fe87",
   124 => x"fe058bc1",
   125 => x"48c087fd",
   126 => x"1e87e6fc",
   127 => x"d4ff1e73",
   128 => x"78ffc348",
   129 => x"1ec04bd3",
   130 => x"c1f0ffc0",
   131 => x"d4fc49c1",
   132 => x"7086c487",
   133 => x"87ca0598",
   134 => x"c348d4ff",
   135 => x"48c178ff",
   136 => x"f1fd87cb",
   137 => x"058bc187",
   138 => x"c087dbff",
   139 => x"87f1fb48",
   140 => x"5c5b5e0e",
   141 => x"4cd4ff0e",
   142 => x"c687dbfd",
   143 => x"e1c01eea",
   144 => x"49c8c1f0",
   145 => x"c487defb",
   146 => x"02a8c186",
   147 => x"eafe87c8",
   148 => x"c148c087",
   149 => x"dafa87e2",
   150 => x"cf497087",
   151 => x"c699ffff",
   152 => x"c802a9ea",
   153 => x"87d3fe87",
   154 => x"cbc148c0",
   155 => x"7cffc387",
   156 => x"fc4bf1c0",
   157 => x"987087f4",
   158 => x"87ebc002",
   159 => x"ffc01ec0",
   160 => x"49fac1f0",
   161 => x"c487defa",
   162 => x"05987086",
   163 => x"ffc387d9",
   164 => x"c3496c7c",
   165 => x"7c7c7cff",
   166 => x"99c0c17c",
   167 => x"c187c402",
   168 => x"c087d548",
   169 => x"c287d148",
   170 => x"87c405ab",
   171 => x"87c848c0",
   172 => x"fe058bc1",
   173 => x"48c087fd",
   174 => x"1e87e4f9",
   175 => x"dcc21e73",
   176 => x"78c148e8",
   177 => x"d0ff4bc7",
   178 => x"fb78c248",
   179 => x"d0ff87c8",
   180 => x"c078c348",
   181 => x"d0e5c01e",
   182 => x"f949c0c1",
   183 => x"86c487c7",
   184 => x"c105a8c1",
   185 => x"abc24b87",
   186 => x"c087c505",
   187 => x"87f9c048",
   188 => x"ff058bc1",
   189 => x"f7fc87d0",
   190 => x"ecdcc287",
   191 => x"05987058",
   192 => x"1ec187cd",
   193 => x"c1f0ffc0",
   194 => x"d8f849d0",
   195 => x"ff86c487",
   196 => x"ffc348d4",
   197 => x"87e0c478",
   198 => x"58f0dcc2",
   199 => x"c248d0ff",
   200 => x"48d4ff78",
   201 => x"c178ffc3",
   202 => x"87f5f748",
   203 => x"5c5b5e0e",
   204 => x"4a710e5d",
   205 => x"ff4dffc3",
   206 => x"7c754cd4",
   207 => x"c448d0ff",
   208 => x"7c7578c3",
   209 => x"ffc01e72",
   210 => x"49d8c1f0",
   211 => x"c487d6f7",
   212 => x"02987086",
   213 => x"48c087c5",
   214 => x"7587f0c0",
   215 => x"7cfec37c",
   216 => x"d41ec0c8",
   217 => x"dcf54966",
   218 => x"7586c487",
   219 => x"757c757c",
   220 => x"e0dad87c",
   221 => x"6c7c754b",
   222 => x"c5059949",
   223 => x"058bc187",
   224 => x"7c7587f3",
   225 => x"c248d0ff",
   226 => x"f648c178",
   227 => x"ff1e87cf",
   228 => x"d0ff4ad4",
   229 => x"78d1c448",
   230 => x"c17affc3",
   231 => x"87f80589",
   232 => x"731e4f26",
   233 => x"c54b711e",
   234 => x"4adfcdee",
   235 => x"c348d4ff",
   236 => x"486878ff",
   237 => x"02a8fec3",
   238 => x"8ac187c5",
   239 => x"7287ed05",
   240 => x"87c5059a",
   241 => x"eac048c0",
   242 => x"029b7387",
   243 => x"66c887cc",
   244 => x"f449731e",
   245 => x"86c487c5",
   246 => x"66c887c6",
   247 => x"87eefe49",
   248 => x"c348d4ff",
   249 => x"737878ff",
   250 => x"87c5059b",
   251 => x"d048d0ff",
   252 => x"f448c178",
   253 => x"731e87eb",
   254 => x"c04a711e",
   255 => x"48d4ff4b",
   256 => x"ff78ffc3",
   257 => x"c3c448d0",
   258 => x"48d4ff78",
   259 => x"7278ffc3",
   260 => x"f0ffc01e",
   261 => x"f449d1c1",
   262 => x"86c487cb",
   263 => x"cd059870",
   264 => x"1ec0c887",
   265 => x"fd4966cc",
   266 => x"86c487f8",
   267 => x"d0ff4b70",
   268 => x"7378c248",
   269 => x"87e9f348",
   270 => x"5c5b5e0e",
   271 => x"1ec00e5d",
   272 => x"c1f0ffc0",
   273 => x"dcf349c9",
   274 => x"c21ed287",
   275 => x"fd49f0dc",
   276 => x"86c887d0",
   277 => x"84c14cc0",
   278 => x"04acb7d2",
   279 => x"dcc287f8",
   280 => x"49bf97f0",
   281 => x"c199c0c3",
   282 => x"c005a9c0",
   283 => x"dcc287e7",
   284 => x"49bf97f7",
   285 => x"dcc231d0",
   286 => x"4abf97f8",
   287 => x"b17232c8",
   288 => x"97f9dcc2",
   289 => x"71b14abf",
   290 => x"ffffcf4c",
   291 => x"84c19cff",
   292 => x"e7c134ca",
   293 => x"f9dcc287",
   294 => x"c149bf97",
   295 => x"c299c631",
   296 => x"bf97fadc",
   297 => x"2ab7c74a",
   298 => x"dcc2b172",
   299 => x"4abf97f5",
   300 => x"c29dcf4d",
   301 => x"bf97f6dc",
   302 => x"ca9ac34a",
   303 => x"f7dcc232",
   304 => x"c24bbf97",
   305 => x"c2b27333",
   306 => x"bf97f8dc",
   307 => x"9bc0c34b",
   308 => x"732bb7c6",
   309 => x"c181c2b2",
   310 => x"70307148",
   311 => x"7548c149",
   312 => x"724d7030",
   313 => x"7184c14c",
   314 => x"b7c0c894",
   315 => x"87cc06ad",
   316 => x"2db734c1",
   317 => x"adb7c0c8",
   318 => x"87f4ff01",
   319 => x"dcf04874",
   320 => x"5b5e0e87",
   321 => x"f80e5d5c",
   322 => x"d6e5c286",
   323 => x"c278c048",
   324 => x"c01ecedd",
   325 => x"87defb49",
   326 => x"987086c4",
   327 => x"c087c505",
   328 => x"87cec948",
   329 => x"7ec14dc0",
   330 => x"bfcbf2c0",
   331 => x"c4dec249",
   332 => x"4bc8714a",
   333 => x"7087f3ec",
   334 => x"87c20598",
   335 => x"f2c07ec0",
   336 => x"c249bfc7",
   337 => x"714ae0de",
   338 => x"ddec4bc8",
   339 => x"05987087",
   340 => x"7ec087c2",
   341 => x"fdc0026e",
   342 => x"d4e4c287",
   343 => x"e5c24dbf",
   344 => x"7ebf9fcc",
   345 => x"ead6c548",
   346 => x"87c705a8",
   347 => x"bfd4e4c2",
   348 => x"6e87ce4d",
   349 => x"d5e9ca48",
   350 => x"87c502a8",
   351 => x"f1c748c0",
   352 => x"ceddc287",
   353 => x"f949751e",
   354 => x"86c487ec",
   355 => x"c5059870",
   356 => x"c748c087",
   357 => x"f2c087dc",
   358 => x"c249bfc7",
   359 => x"714ae0de",
   360 => x"c5eb4bc8",
   361 => x"05987087",
   362 => x"e5c287c8",
   363 => x"78c148d6",
   364 => x"f2c087da",
   365 => x"c249bfcb",
   366 => x"714ac4de",
   367 => x"e9ea4bc8",
   368 => x"02987087",
   369 => x"c087c5c0",
   370 => x"87e6c648",
   371 => x"97cce5c2",
   372 => x"d5c149bf",
   373 => x"cdc005a9",
   374 => x"cde5c287",
   375 => x"c249bf97",
   376 => x"c002a9ea",
   377 => x"48c087c5",
   378 => x"c287c7c6",
   379 => x"bf97cedd",
   380 => x"e9c3487e",
   381 => x"cec002a8",
   382 => x"c3486e87",
   383 => x"c002a8eb",
   384 => x"48c087c5",
   385 => x"c287ebc5",
   386 => x"bf97d9dd",
   387 => x"c0059949",
   388 => x"ddc287cc",
   389 => x"49bf97da",
   390 => x"c002a9c2",
   391 => x"48c087c5",
   392 => x"c287cfc5",
   393 => x"bf97dbdd",
   394 => x"d2e5c248",
   395 => x"484c7058",
   396 => x"e5c288c1",
   397 => x"ddc258d6",
   398 => x"49bf97dc",
   399 => x"ddc28175",
   400 => x"4abf97dd",
   401 => x"a17232c8",
   402 => x"e3e9c27e",
   403 => x"c2786e48",
   404 => x"bf97dedd",
   405 => x"58a6c848",
   406 => x"bfd6e5c2",
   407 => x"87d4c202",
   408 => x"bfc7f2c0",
   409 => x"e0dec249",
   410 => x"4bc8714a",
   411 => x"7087fbe7",
   412 => x"c5c00298",
   413 => x"c348c087",
   414 => x"e5c287f8",
   415 => x"c24cbfce",
   416 => x"c25cf7e9",
   417 => x"bf97f3dd",
   418 => x"c231c849",
   419 => x"bf97f2dd",
   420 => x"c249a14a",
   421 => x"bf97f4dd",
   422 => x"7232d04a",
   423 => x"ddc249a1",
   424 => x"4abf97f5",
   425 => x"a17232d8",
   426 => x"9166c449",
   427 => x"bfe3e9c2",
   428 => x"ebe9c281",
   429 => x"fbddc259",
   430 => x"c84abf97",
   431 => x"faddc232",
   432 => x"a24bbf97",
   433 => x"fcddc24a",
   434 => x"d04bbf97",
   435 => x"4aa27333",
   436 => x"97fdddc2",
   437 => x"9bcf4bbf",
   438 => x"a27333d8",
   439 => x"efe9c24a",
   440 => x"ebe9c25a",
   441 => x"8ac24abf",
   442 => x"e9c29274",
   443 => x"a17248ef",
   444 => x"87cac178",
   445 => x"97e0ddc2",
   446 => x"31c849bf",
   447 => x"97dfddc2",
   448 => x"49a14abf",
   449 => x"59dee5c2",
   450 => x"bfdae5c2",
   451 => x"c731c549",
   452 => x"29c981ff",
   453 => x"59f7e9c2",
   454 => x"97e5ddc2",
   455 => x"32c84abf",
   456 => x"97e4ddc2",
   457 => x"4aa24bbf",
   458 => x"6e9266c4",
   459 => x"f3e9c282",
   460 => x"ebe9c25a",
   461 => x"c278c048",
   462 => x"7248e7e9",
   463 => x"e9c278a1",
   464 => x"e9c248f7",
   465 => x"c278bfeb",
   466 => x"c248fbe9",
   467 => x"78bfefe9",
   468 => x"bfd6e5c2",
   469 => x"87c9c002",
   470 => x"30c44874",
   471 => x"c9c07e70",
   472 => x"f3e9c287",
   473 => x"30c448bf",
   474 => x"e5c27e70",
   475 => x"786e48da",
   476 => x"8ef848c1",
   477 => x"4c264d26",
   478 => x"4f264b26",
   479 => x"5c5b5e0e",
   480 => x"4a710e5d",
   481 => x"bfd6e5c2",
   482 => x"7287cb02",
   483 => x"722bc74b",
   484 => x"9cffc14c",
   485 => x"4b7287c9",
   486 => x"4c722bc8",
   487 => x"c29cffc3",
   488 => x"83bfe3e9",
   489 => x"bfc3f2c0",
   490 => x"87d902ab",
   491 => x"5bc7f2c0",
   492 => x"1eceddc2",
   493 => x"fdf04973",
   494 => x"7086c487",
   495 => x"87c50598",
   496 => x"e6c048c0",
   497 => x"d6e5c287",
   498 => x"87d202bf",
   499 => x"91c44974",
   500 => x"81ceddc2",
   501 => x"ffcf4d69",
   502 => x"9dffffff",
   503 => x"497487cb",
   504 => x"ddc291c2",
   505 => x"699f81ce",
   506 => x"fe48754d",
   507 => x"5e0e87c6",
   508 => x"0e5d5c5b",
   509 => x"c04d711e",
   510 => x"ca49c11e",
   511 => x"86c487ee",
   512 => x"029c4c70",
   513 => x"c287c0c1",
   514 => x"754adee5",
   515 => x"87ffe049",
   516 => x"c0029870",
   517 => x"4a7487f1",
   518 => x"4bcb4975",
   519 => x"7087e5e1",
   520 => x"e2c00298",
   521 => x"741ec087",
   522 => x"87c7029c",
   523 => x"c048a6c4",
   524 => x"c487c578",
   525 => x"78c148a6",
   526 => x"c94966c4",
   527 => x"86c487ee",
   528 => x"059c4c70",
   529 => x"7487c0ff",
   530 => x"e7fc2648",
   531 => x"5b5e0e87",
   532 => x"1e0e5d5c",
   533 => x"059b4b71",
   534 => x"48c087c5",
   535 => x"c887e5c1",
   536 => x"7dc04da3",
   537 => x"c70266d4",
   538 => x"9766d487",
   539 => x"87c505bf",
   540 => x"cfc148c0",
   541 => x"4966d487",
   542 => x"7087f3fd",
   543 => x"c1029c4c",
   544 => x"a4dc87c0",
   545 => x"da7d6949",
   546 => x"a3c449a4",
   547 => x"7a699f4a",
   548 => x"bfd6e5c2",
   549 => x"d487d202",
   550 => x"699f49a4",
   551 => x"ffffc049",
   552 => x"d0487199",
   553 => x"c27e7030",
   554 => x"6e7ec087",
   555 => x"806a4849",
   556 => x"7bc07a70",
   557 => x"6a49a3cc",
   558 => x"49a3d079",
   559 => x"487479c0",
   560 => x"48c087c2",
   561 => x"87ecfa26",
   562 => x"5c5b5e0e",
   563 => x"4c710e5d",
   564 => x"48c3f2c0",
   565 => x"9c7478ff",
   566 => x"87cac102",
   567 => x"6949a4c8",
   568 => x"87c2c102",
   569 => x"6c4a66d0",
   570 => x"a6d48249",
   571 => x"4d66d05a",
   572 => x"d2e5c2b9",
   573 => x"baff4abf",
   574 => x"99719972",
   575 => x"87e4c002",
   576 => x"6b4ba4c4",
   577 => x"87f4f949",
   578 => x"e5c27b70",
   579 => x"6c49bfce",
   580 => x"757c7181",
   581 => x"d2e5c2b9",
   582 => x"baff4abf",
   583 => x"99719972",
   584 => x"87dcff05",
   585 => x"cbf97c75",
   586 => x"1e731e87",
   587 => x"029b4b71",
   588 => x"a3c887c7",
   589 => x"c5056949",
   590 => x"c048c087",
   591 => x"e9c287eb",
   592 => x"c44abfe7",
   593 => x"496949a3",
   594 => x"e5c289c2",
   595 => x"7191bfce",
   596 => x"e5c24aa2",
   597 => x"6b49bfd2",
   598 => x"4aa27199",
   599 => x"721e66c8",
   600 => x"87d2ea49",
   601 => x"497086c4",
   602 => x"87ccf848",
   603 => x"711e731e",
   604 => x"c7029b4b",
   605 => x"49a3c887",
   606 => x"87c50569",
   607 => x"ebc048c0",
   608 => x"e7e9c287",
   609 => x"a3c44abf",
   610 => x"c2496949",
   611 => x"cee5c289",
   612 => x"a27191bf",
   613 => x"d2e5c24a",
   614 => x"996b49bf",
   615 => x"c84aa271",
   616 => x"49721e66",
   617 => x"c487c5e6",
   618 => x"48497086",
   619 => x"0e87c9f7",
   620 => x"5d5c5b5e",
   621 => x"4b711e0e",
   622 => x"c94c66d4",
   623 => x"029b732c",
   624 => x"c887cfc1",
   625 => x"026949a3",
   626 => x"d087c7c1",
   627 => x"66d44da3",
   628 => x"d2e5c27d",
   629 => x"b9ff49bf",
   630 => x"7e994a6b",
   631 => x"cd03ac71",
   632 => x"7d7bc087",
   633 => x"c44aa3cc",
   634 => x"796a49a3",
   635 => x"8c7287c2",
   636 => x"dd029c74",
   637 => x"731e4987",
   638 => x"87ccfb49",
   639 => x"66d486c4",
   640 => x"99ffc749",
   641 => x"c287cb02",
   642 => x"731ecedd",
   643 => x"87d9fc49",
   644 => x"f52686c4",
   645 => x"731e87de",
   646 => x"9b4b711e",
   647 => x"87e4c002",
   648 => x"5bfbe9c2",
   649 => x"8ac24a73",
   650 => x"bfcee5c2",
   651 => x"e9c29249",
   652 => x"7248bfe7",
   653 => x"ffe9c280",
   654 => x"c4487158",
   655 => x"dee5c230",
   656 => x"87edc058",
   657 => x"48f7e9c2",
   658 => x"bfebe9c2",
   659 => x"fbe9c278",
   660 => x"efe9c248",
   661 => x"e5c278bf",
   662 => x"c902bfd6",
   663 => x"cee5c287",
   664 => x"31c449bf",
   665 => x"e9c287c7",
   666 => x"c449bff3",
   667 => x"dee5c231",
   668 => x"87c4f459",
   669 => x"5c5b5e0e",
   670 => x"c04a710e",
   671 => x"029a724b",
   672 => x"da87e1c0",
   673 => x"699f49a2",
   674 => x"d6e5c24b",
   675 => x"87cf02bf",
   676 => x"9f49a2d4",
   677 => x"c04c4969",
   678 => x"d09cffff",
   679 => x"c087c234",
   680 => x"b349744c",
   681 => x"edfd4973",
   682 => x"87caf387",
   683 => x"5c5b5e0e",
   684 => x"86f40e5d",
   685 => x"7ec04a71",
   686 => x"d8029a72",
   687 => x"caddc287",
   688 => x"c278c048",
   689 => x"c248c2dd",
   690 => x"78bffbe9",
   691 => x"48c6ddc2",
   692 => x"bff7e9c2",
   693 => x"ebe5c278",
   694 => x"c250c048",
   695 => x"49bfdae5",
   696 => x"bfcaddc2",
   697 => x"03aa714a",
   698 => x"7287ffc3",
   699 => x"0599cf49",
   700 => x"c287e0c0",
   701 => x"c21ecedd",
   702 => x"49bfc2dd",
   703 => x"48c2ddc2",
   704 => x"7178a1c1",
   705 => x"c487efe3",
   706 => x"fff1c086",
   707 => x"ceddc248",
   708 => x"c087cc78",
   709 => x"48bffff1",
   710 => x"c080e0c0",
   711 => x"c258c3f2",
   712 => x"48bfcadd",
   713 => x"ddc280c1",
   714 => x"7f2758ce",
   715 => x"bf00000c",
   716 => x"9d4dbf97",
   717 => x"87e2c202",
   718 => x"02ade5c3",
   719 => x"c087dbc2",
   720 => x"4bbffff1",
   721 => x"1149a3cb",
   722 => x"05accf4c",
   723 => x"7587d2c1",
   724 => x"c199df49",
   725 => x"c291cd89",
   726 => x"c181dee5",
   727 => x"51124aa3",
   728 => x"124aa3c3",
   729 => x"4aa3c551",
   730 => x"a3c75112",
   731 => x"c951124a",
   732 => x"51124aa3",
   733 => x"124aa3ce",
   734 => x"4aa3d051",
   735 => x"a3d25112",
   736 => x"d451124a",
   737 => x"51124aa3",
   738 => x"124aa3d6",
   739 => x"4aa3d851",
   740 => x"a3dc5112",
   741 => x"de51124a",
   742 => x"51124aa3",
   743 => x"f9c07ec1",
   744 => x"c8497487",
   745 => x"eac00599",
   746 => x"d0497487",
   747 => x"87d00599",
   748 => x"c00266dc",
   749 => x"497387ca",
   750 => x"700f66dc",
   751 => x"87d30298",
   752 => x"c6c0056e",
   753 => x"dee5c287",
   754 => x"c050c048",
   755 => x"48bffff1",
   756 => x"c287e7c2",
   757 => x"c048ebe5",
   758 => x"e5c27e50",
   759 => x"c249bfda",
   760 => x"4abfcadd",
   761 => x"fc04aa71",
   762 => x"e9c287c1",
   763 => x"c005bffb",
   764 => x"e5c287c8",
   765 => x"c102bfd6",
   766 => x"f2c087fe",
   767 => x"78ff48c3",
   768 => x"bfc6ddc2",
   769 => x"87f4ed49",
   770 => x"ddc24970",
   771 => x"a6c459ca",
   772 => x"c6ddc248",
   773 => x"e5c278bf",
   774 => x"c002bfd6",
   775 => x"66c487d8",
   776 => x"ffffcf49",
   777 => x"a999f8ff",
   778 => x"87c5c002",
   779 => x"e1c04dc0",
   780 => x"c04dc187",
   781 => x"66c487dc",
   782 => x"f8ffcf49",
   783 => x"c002a999",
   784 => x"a6c887c8",
   785 => x"c078c048",
   786 => x"a6c887c5",
   787 => x"c878c148",
   788 => x"9d754d66",
   789 => x"87e0c005",
   790 => x"c24966c4",
   791 => x"cee5c289",
   792 => x"c2914abf",
   793 => x"4abfe7e9",
   794 => x"48c2ddc2",
   795 => x"c278a172",
   796 => x"c048cadd",
   797 => x"87e3f978",
   798 => x"8ef448c0",
   799 => x"0087f5eb",
   800 => x"ff000000",
   801 => x"8fffffff",
   802 => x"9800000c",
   803 => x"4600000c",
   804 => x"32335441",
   805 => x"00202020",
   806 => x"31544146",
   807 => x"20202036",
   808 => x"d4ff1e00",
   809 => x"78ffc348",
   810 => x"4f264868",
   811 => x"48d4ff1e",
   812 => x"ff78ffc3",
   813 => x"e1c848d0",
   814 => x"48d4ff78",
   815 => x"e9c278d4",
   816 => x"d4ff48ff",
   817 => x"4f2650bf",
   818 => x"48d0ff1e",
   819 => x"2678e0c0",
   820 => x"ccff1e4f",
   821 => x"99497087",
   822 => x"c087c602",
   823 => x"f105a9fb",
   824 => x"26487187",
   825 => x"5b5e0e4f",
   826 => x"4b710e5c",
   827 => x"f0fe4cc0",
   828 => x"99497087",
   829 => x"87f9c002",
   830 => x"02a9ecc0",
   831 => x"c087f2c0",
   832 => x"c002a9fb",
   833 => x"66cc87eb",
   834 => x"c703acb7",
   835 => x"0266d087",
   836 => x"537187c2",
   837 => x"c2029971",
   838 => x"fe84c187",
   839 => x"497087c3",
   840 => x"87cd0299",
   841 => x"02a9ecc0",
   842 => x"fbc087c7",
   843 => x"d5ff05a9",
   844 => x"0266d087",
   845 => x"97c087c3",
   846 => x"a9ecc07b",
   847 => x"7487c405",
   848 => x"7487c54a",
   849 => x"8a0ac04a",
   850 => x"87c24872",
   851 => x"4c264d26",
   852 => x"4f264b26",
   853 => x"87c9fd1e",
   854 => x"f0c04970",
   855 => x"ca04a9b7",
   856 => x"b7f9c087",
   857 => x"87c301a9",
   858 => x"c189f0c0",
   859 => x"04a9b7c1",
   860 => x"dac187ca",
   861 => x"c301a9b7",
   862 => x"89f7c087",
   863 => x"4f264871",
   864 => x"5c5b5e0e",
   865 => x"ff4a710e",
   866 => x"49724cd4",
   867 => x"7087eac0",
   868 => x"c2029b4b",
   869 => x"ff8bc187",
   870 => x"c5c848d0",
   871 => x"7cd5c178",
   872 => x"31c64973",
   873 => x"97d2dbc2",
   874 => x"71484abf",
   875 => x"ff7c70b0",
   876 => x"78c448d0",
   877 => x"d5fe4873",
   878 => x"5b5e0e87",
   879 => x"f80e5d5c",
   880 => x"c04c7186",
   881 => x"87e4fb7e",
   882 => x"f9c04bc0",
   883 => x"49bf97e6",
   884 => x"cf04a9c0",
   885 => x"87f9fb87",
   886 => x"f9c083c1",
   887 => x"49bf97e6",
   888 => x"87f106ab",
   889 => x"97e6f9c0",
   890 => x"87cf02bf",
   891 => x"7087f2fa",
   892 => x"c6029949",
   893 => x"a9ecc087",
   894 => x"c087f105",
   895 => x"87e1fa4b",
   896 => x"dcfa4d70",
   897 => x"58a6c887",
   898 => x"7087d6fa",
   899 => x"c883c14a",
   900 => x"699749a4",
   901 => x"c702ad49",
   902 => x"adffc087",
   903 => x"87e7c005",
   904 => x"9749a4c9",
   905 => x"66c44969",
   906 => x"87c702a9",
   907 => x"a8ffc048",
   908 => x"ca87d405",
   909 => x"699749a4",
   910 => x"c602aa49",
   911 => x"aaffc087",
   912 => x"c187c405",
   913 => x"c087d07e",
   914 => x"c602adec",
   915 => x"adfbc087",
   916 => x"c087c405",
   917 => x"6e7ec14b",
   918 => x"87e1fe02",
   919 => x"7387e9f9",
   920 => x"fb8ef848",
   921 => x"0e0087e6",
   922 => x"5d5c5b5e",
   923 => x"4b711e0e",
   924 => x"ab4d4cc0",
   925 => x"87e8c004",
   926 => x"1ef9f6c0",
   927 => x"c4029d75",
   928 => x"c24ac087",
   929 => x"724ac187",
   930 => x"87e0f049",
   931 => x"7e7086c4",
   932 => x"056e84c1",
   933 => x"4c7387c2",
   934 => x"ac7385c1",
   935 => x"87d8ff06",
   936 => x"2626486e",
   937 => x"264c264d",
   938 => x"0e4f264b",
   939 => x"5d5c5b5e",
   940 => x"4c711e0e",
   941 => x"c291de49",
   942 => x"714dd9ea",
   943 => x"026d9785",
   944 => x"c287ddc1",
   945 => x"4abfc4ea",
   946 => x"49728274",
   947 => x"7087d8fe",
   948 => x"c0026e7e",
   949 => x"eac287f3",
   950 => x"4a6e4bcc",
   951 => x"c7ff49cb",
   952 => x"4b7487c6",
   953 => x"ddc193cb",
   954 => x"83c483fa",
   955 => x"7be4fcc0",
   956 => x"c3c14974",
   957 => x"7b7587f3",
   958 => x"97d8eac2",
   959 => x"c21e49bf",
   960 => x"c149ccea",
   961 => x"c487cdde",
   962 => x"c1497486",
   963 => x"c087dac3",
   964 => x"f9c4c149",
   965 => x"c0eac287",
   966 => x"c178c048",
   967 => x"87cbdd49",
   968 => x"87fffd26",
   969 => x"64616f4c",
   970 => x"2e676e69",
   971 => x"0e002e2e",
   972 => x"0e5c5b5e",
   973 => x"c24a4b71",
   974 => x"82bfc4ea",
   975 => x"e6fc4972",
   976 => x"9c4c7087",
   977 => x"4987c402",
   978 => x"c287e9ec",
   979 => x"c048c4ea",
   980 => x"dc49c178",
   981 => x"ccfd87d5",
   982 => x"5b5e0e87",
   983 => x"f40e5d5c",
   984 => x"ceddc286",
   985 => x"c44cc04d",
   986 => x"78c048a6",
   987 => x"bfc4eac2",
   988 => x"06a9c049",
   989 => x"c287c1c1",
   990 => x"9848cedd",
   991 => x"87f8c002",
   992 => x"1ef9f6c0",
   993 => x"c70266c8",
   994 => x"48a6c487",
   995 => x"87c578c0",
   996 => x"c148a6c4",
   997 => x"4966c478",
   998 => x"c487d1ec",
   999 => x"c14d7086",
  1000 => x"4866c484",
  1001 => x"a6c880c1",
  1002 => x"c4eac258",
  1003 => x"03ac49bf",
  1004 => x"9d7587c6",
  1005 => x"87c8ff05",
  1006 => x"9d754cc0",
  1007 => x"87e0c302",
  1008 => x"1ef9f6c0",
  1009 => x"c70266c8",
  1010 => x"48a6cc87",
  1011 => x"87c578c0",
  1012 => x"c148a6cc",
  1013 => x"4966cc78",
  1014 => x"c487d1eb",
  1015 => x"6e7e7086",
  1016 => x"87e9c202",
  1017 => x"81cb496e",
  1018 => x"d0496997",
  1019 => x"d6c10299",
  1020 => x"effcc087",
  1021 => x"cb49744a",
  1022 => x"faddc191",
  1023 => x"c8797281",
  1024 => x"51ffc381",
  1025 => x"91de4974",
  1026 => x"4dd9eac2",
  1027 => x"c1c28571",
  1028 => x"a5c17d97",
  1029 => x"51e0c049",
  1030 => x"97dee5c2",
  1031 => x"87d202bf",
  1032 => x"a5c284c1",
  1033 => x"dee5c24b",
  1034 => x"ff49db4a",
  1035 => x"c187f9c1",
  1036 => x"a5cd87db",
  1037 => x"c151c049",
  1038 => x"4ba5c284",
  1039 => x"49cb4a6e",
  1040 => x"87e4c1ff",
  1041 => x"c087c6c1",
  1042 => x"744aebfa",
  1043 => x"c191cb49",
  1044 => x"7281fadd",
  1045 => x"dee5c279",
  1046 => x"d802bf97",
  1047 => x"de497487",
  1048 => x"c284c191",
  1049 => x"714bd9ea",
  1050 => x"dee5c283",
  1051 => x"ff49dd4a",
  1052 => x"d887f5c0",
  1053 => x"de4b7487",
  1054 => x"d9eac293",
  1055 => x"49a3cb83",
  1056 => x"84c151c0",
  1057 => x"cb4a6e73",
  1058 => x"dbc0ff49",
  1059 => x"4866c487",
  1060 => x"a6c880c1",
  1061 => x"03acc758",
  1062 => x"6e87c5c0",
  1063 => x"87e0fc05",
  1064 => x"8ef44874",
  1065 => x"1e87fcf7",
  1066 => x"4b711e73",
  1067 => x"c191cb49",
  1068 => x"c881fadd",
  1069 => x"dbc24aa1",
  1070 => x"501248d2",
  1071 => x"c04aa1c9",
  1072 => x"1248e6f9",
  1073 => x"c281ca50",
  1074 => x"1148d8ea",
  1075 => x"d8eac250",
  1076 => x"1e49bf97",
  1077 => x"d6c149c0",
  1078 => x"eac287fa",
  1079 => x"78de48c0",
  1080 => x"c6d649c1",
  1081 => x"fef62687",
  1082 => x"4a711e87",
  1083 => x"c191cb49",
  1084 => x"c881fadd",
  1085 => x"c2481181",
  1086 => x"c258c4ea",
  1087 => x"c048c4ea",
  1088 => x"d549c178",
  1089 => x"4f2687e5",
  1090 => x"c049c01e",
  1091 => x"2687fffc",
  1092 => x"99711e4f",
  1093 => x"c187d202",
  1094 => x"c048cfdf",
  1095 => x"c180f750",
  1096 => x"c140e9c3",
  1097 => x"ce78f3dd",
  1098 => x"cbdfc187",
  1099 => x"ecddc148",
  1100 => x"c180fc78",
  1101 => x"2678c8c4",
  1102 => x"5b5e0e4f",
  1103 => x"4c710e5c",
  1104 => x"c192cb4a",
  1105 => x"c882fadd",
  1106 => x"a2c949a2",
  1107 => x"4b6b974b",
  1108 => x"4969971e",
  1109 => x"1282ca1e",
  1110 => x"fae7c049",
  1111 => x"d449c087",
  1112 => x"497487c9",
  1113 => x"87c1fac0",
  1114 => x"f8f48ef8",
  1115 => x"1e731e87",
  1116 => x"ff494b71",
  1117 => x"497387c3",
  1118 => x"f487fefe",
  1119 => x"731e87e9",
  1120 => x"c64b711e",
  1121 => x"db024aa3",
  1122 => x"028ac187",
  1123 => x"028a87d6",
  1124 => x"8a87dac1",
  1125 => x"87fcc002",
  1126 => x"e1c0028a",
  1127 => x"cb028a87",
  1128 => x"87dbc187",
  1129 => x"c0fd49c7",
  1130 => x"87dec187",
  1131 => x"bfc4eac2",
  1132 => x"87cbc102",
  1133 => x"c288c148",
  1134 => x"c158c8ea",
  1135 => x"eac287c1",
  1136 => x"c002bfc8",
  1137 => x"eac287f9",
  1138 => x"c148bfc4",
  1139 => x"c8eac280",
  1140 => x"87ebc058",
  1141 => x"bfc4eac2",
  1142 => x"c289c649",
  1143 => x"c059c8ea",
  1144 => x"da03a9b7",
  1145 => x"c4eac287",
  1146 => x"d278c048",
  1147 => x"c8eac287",
  1148 => x"87cb02bf",
  1149 => x"bfc4eac2",
  1150 => x"c280c648",
  1151 => x"c058c8ea",
  1152 => x"87e7d149",
  1153 => x"f7c04973",
  1154 => x"daf287df",
  1155 => x"5b5e0e87",
  1156 => x"4c710e5c",
  1157 => x"741e66cc",
  1158 => x"c193cb4b",
  1159 => x"c483fadd",
  1160 => x"496a4aa3",
  1161 => x"87d0fafe",
  1162 => x"7be7c2c1",
  1163 => x"d449a3c8",
  1164 => x"a3c95166",
  1165 => x"5166d849",
  1166 => x"dc49a3ca",
  1167 => x"f1265166",
  1168 => x"5e0e87e3",
  1169 => x"0e5d5c5b",
  1170 => x"d886d0ff",
  1171 => x"a6c459a6",
  1172 => x"c478c048",
  1173 => x"66c4c180",
  1174 => x"c180c478",
  1175 => x"c180c478",
  1176 => x"c8eac278",
  1177 => x"c278c148",
  1178 => x"48bfc0ea",
  1179 => x"cb05a8de",
  1180 => x"87e5f387",
  1181 => x"a6c84970",
  1182 => x"87f8ce59",
  1183 => x"e987ede8",
  1184 => x"dce887cf",
  1185 => x"c04c7087",
  1186 => x"c102acfb",
  1187 => x"66d487d0",
  1188 => x"87c2c105",
  1189 => x"c11e1ec0",
  1190 => x"eddfc11e",
  1191 => x"fd49c01e",
  1192 => x"d0c187eb",
  1193 => x"82c44a66",
  1194 => x"81c7496a",
  1195 => x"1ec15174",
  1196 => x"496a1ed8",
  1197 => x"ece881c8",
  1198 => x"c186d887",
  1199 => x"c04866c4",
  1200 => x"87c701a8",
  1201 => x"c148a6c4",
  1202 => x"c187ce78",
  1203 => x"c14866c4",
  1204 => x"58a6cc88",
  1205 => x"f8e787c3",
  1206 => x"48a6cc87",
  1207 => x"9c7478c2",
  1208 => x"87cccd02",
  1209 => x"c14866c4",
  1210 => x"03a866c8",
  1211 => x"d887c1cd",
  1212 => x"78c048a6",
  1213 => x"7087eae6",
  1214 => x"acd0c14c",
  1215 => x"87d6c205",
  1216 => x"e97e66d8",
  1217 => x"497087ce",
  1218 => x"e659a6dc",
  1219 => x"4c7087d3",
  1220 => x"05acecc0",
  1221 => x"c487eac1",
  1222 => x"91cb4966",
  1223 => x"8166c0c1",
  1224 => x"6a4aa1c4",
  1225 => x"4aa1c84d",
  1226 => x"c15266d8",
  1227 => x"e579e9c3",
  1228 => x"4c7087ef",
  1229 => x"87d8029c",
  1230 => x"02acfbc0",
  1231 => x"557487d2",
  1232 => x"7087dee5",
  1233 => x"c7029c4c",
  1234 => x"acfbc087",
  1235 => x"87eeff05",
  1236 => x"c255e0c0",
  1237 => x"97c055c1",
  1238 => x"4966d47d",
  1239 => x"db05a96e",
  1240 => x"4866c487",
  1241 => x"04a866c8",
  1242 => x"66c487ca",
  1243 => x"c880c148",
  1244 => x"87c858a6",
  1245 => x"c14866c8",
  1246 => x"58a6cc88",
  1247 => x"7087e2e4",
  1248 => x"acd0c14c",
  1249 => x"d087c805",
  1250 => x"80c14866",
  1251 => x"c158a6d4",
  1252 => x"fd02acd0",
  1253 => x"a6dc87ea",
  1254 => x"7866d448",
  1255 => x"dc4866d8",
  1256 => x"c905a866",
  1257 => x"e0c087dc",
  1258 => x"f0c048a6",
  1259 => x"cc80c478",
  1260 => x"80c47866",
  1261 => x"747e78c0",
  1262 => x"88fbc048",
  1263 => x"58a6f0c0",
  1264 => x"c8029870",
  1265 => x"cb4887d7",
  1266 => x"a6f0c088",
  1267 => x"02987058",
  1268 => x"4887e9c0",
  1269 => x"f0c088c9",
  1270 => x"987058a6",
  1271 => x"87e1c302",
  1272 => x"c088c448",
  1273 => x"7058a6f0",
  1274 => x"87de0298",
  1275 => x"c088c148",
  1276 => x"7058a6f0",
  1277 => x"c8c30298",
  1278 => x"87dbc787",
  1279 => x"48a6e0c0",
  1280 => x"66cc78c0",
  1281 => x"d080c148",
  1282 => x"d4e258a6",
  1283 => x"c04c7087",
  1284 => x"d502acec",
  1285 => x"66e0c087",
  1286 => x"c087c602",
  1287 => x"c95ca6e4",
  1288 => x"c0487487",
  1289 => x"e8c088f0",
  1290 => x"ecc058a6",
  1291 => x"87cc02ac",
  1292 => x"7087eee1",
  1293 => x"acecc04c",
  1294 => x"87f4ff05",
  1295 => x"1e66e0c0",
  1296 => x"1e4966d4",
  1297 => x"1e66ecc0",
  1298 => x"1eeddfc1",
  1299 => x"f64966d4",
  1300 => x"1ec087fb",
  1301 => x"66dc1eca",
  1302 => x"c191cb49",
  1303 => x"d88166d8",
  1304 => x"a1c448a6",
  1305 => x"bf66d878",
  1306 => x"87f9e149",
  1307 => x"b7c086d8",
  1308 => x"c7c106a8",
  1309 => x"de1ec187",
  1310 => x"bf66c81e",
  1311 => x"87e5e149",
  1312 => x"497086c8",
  1313 => x"8808c048",
  1314 => x"58a6e4c0",
  1315 => x"06a8b7c0",
  1316 => x"c087e9c0",
  1317 => x"dd4866e0",
  1318 => x"df03a8b7",
  1319 => x"49bf6e87",
  1320 => x"8166e0c0",
  1321 => x"6651e0c0",
  1322 => x"6e81c149",
  1323 => x"c1c281bf",
  1324 => x"66e0c051",
  1325 => x"6e81c249",
  1326 => x"51c081bf",
  1327 => x"dcc47ec1",
  1328 => x"87d0e287",
  1329 => x"58a6e4c0",
  1330 => x"c087c9e2",
  1331 => x"c058a6e8",
  1332 => x"c005a8ec",
  1333 => x"e4c087cb",
  1334 => x"e0c048a6",
  1335 => x"c4c07866",
  1336 => x"fcdeff87",
  1337 => x"4966c487",
  1338 => x"c0c191cb",
  1339 => x"80714866",
  1340 => x"4a6e7e70",
  1341 => x"496e82c8",
  1342 => x"e0c081ca",
  1343 => x"e4c05166",
  1344 => x"81c14966",
  1345 => x"8966e0c0",
  1346 => x"307148c1",
  1347 => x"89c14970",
  1348 => x"c27a9771",
  1349 => x"49bff5ed",
  1350 => x"2966e0c0",
  1351 => x"484a6a97",
  1352 => x"f0c09871",
  1353 => x"496e58a6",
  1354 => x"4d6981c4",
  1355 => x"d84866dc",
  1356 => x"c002a866",
  1357 => x"a6d887c8",
  1358 => x"c078c048",
  1359 => x"a6d887c5",
  1360 => x"d878c148",
  1361 => x"e0c01e66",
  1362 => x"ff49751e",
  1363 => x"c887d6de",
  1364 => x"c04c7086",
  1365 => x"c106acb7",
  1366 => x"857487d4",
  1367 => x"7449e0c0",
  1368 => x"c14b7589",
  1369 => x"714ae8d9",
  1370 => x"87fcecfe",
  1371 => x"e8c085c2",
  1372 => x"80c14866",
  1373 => x"58a6ecc0",
  1374 => x"4966ecc0",
  1375 => x"a97081c1",
  1376 => x"87c8c002",
  1377 => x"c048a6d8",
  1378 => x"87c5c078",
  1379 => x"c148a6d8",
  1380 => x"1e66d878",
  1381 => x"c049a4c2",
  1382 => x"887148e0",
  1383 => x"751e4970",
  1384 => x"c0ddff49",
  1385 => x"c086c887",
  1386 => x"ff01a8b7",
  1387 => x"e8c087c0",
  1388 => x"d1c00266",
  1389 => x"c9496e87",
  1390 => x"66e8c081",
  1391 => x"c1486e51",
  1392 => x"c078f9c4",
  1393 => x"496e87cc",
  1394 => x"51c281c9",
  1395 => x"c5c1486e",
  1396 => x"7ec178ed",
  1397 => x"ff87c6c0",
  1398 => x"7087f6db",
  1399 => x"c0026e4c",
  1400 => x"66c487f5",
  1401 => x"a866c848",
  1402 => x"87cbc004",
  1403 => x"c14866c4",
  1404 => x"58a6c880",
  1405 => x"c887e0c0",
  1406 => x"88c14866",
  1407 => x"c058a6cc",
  1408 => x"c6c187d5",
  1409 => x"c8c005ac",
  1410 => x"4866cc87",
  1411 => x"a6d080c1",
  1412 => x"fcdaff58",
  1413 => x"d04c7087",
  1414 => x"80c14866",
  1415 => x"7458a6d4",
  1416 => x"cbc0029c",
  1417 => x"4866c487",
  1418 => x"a866c8c1",
  1419 => x"87fff204",
  1420 => x"87d4daff",
  1421 => x"c74866c4",
  1422 => x"e5c003a8",
  1423 => x"c8eac287",
  1424 => x"c478c048",
  1425 => x"91cb4966",
  1426 => x"8166c0c1",
  1427 => x"6a4aa1c4",
  1428 => x"7952c04a",
  1429 => x"c14866c4",
  1430 => x"58a6c880",
  1431 => x"ff04a8c7",
  1432 => x"d0ff87db",
  1433 => x"87fbe08e",
  1434 => x"1e00203a",
  1435 => x"4b711e73",
  1436 => x"87c6029b",
  1437 => x"48c4eac2",
  1438 => x"1ec778c0",
  1439 => x"bfc4eac2",
  1440 => x"ddc11e49",
  1441 => x"eac21efa",
  1442 => x"ee49bfc0",
  1443 => x"86cc87f4",
  1444 => x"bfc0eac2",
  1445 => x"87f9e949",
  1446 => x"c8029b73",
  1447 => x"faddc187",
  1448 => x"d6e6c049",
  1449 => x"fedfff87",
  1450 => x"1e731e87",
  1451 => x"dbc24bc0",
  1452 => x"50c048d2",
  1453 => x"bfdddfc1",
  1454 => x"eafbc049",
  1455 => x"05987087",
  1456 => x"dbc187c4",
  1457 => x"48734bcc",
  1458 => x"87dbdfff",
  1459 => x"204d4f52",
  1460 => x"64616f6c",
  1461 => x"20676e69",
  1462 => x"6c696166",
  1463 => x"1e006465",
  1464 => x"c187e9c7",
  1465 => x"87c3fe49",
  1466 => x"87cfeffe",
  1467 => x"cd029870",
  1468 => x"ccf8fe87",
  1469 => x"02987087",
  1470 => x"4ac187c4",
  1471 => x"4ac087c2",
  1472 => x"ce059a72",
  1473 => x"c11ec087",
  1474 => x"c049f3dc",
  1475 => x"c487fbf0",
  1476 => x"c087fe86",
  1477 => x"c087e5ff",
  1478 => x"fedcc11e",
  1479 => x"e9f0c049",
  1480 => x"fe1ec087",
  1481 => x"497087c3",
  1482 => x"87def0c0",
  1483 => x"f887dcc3",
  1484 => x"534f268e",
  1485 => x"61662044",
  1486 => x"64656c69",
  1487 => x"6f42002e",
  1488 => x"6e69746f",
  1489 => x"2e2e2e67",
  1490 => x"e8c01e00",
  1491 => x"f3c087c9",
  1492 => x"87f687ee",
  1493 => x"c21e4f26",
  1494 => x"c048c4ea",
  1495 => x"c0eac278",
  1496 => x"fd78c048",
  1497 => x"87e187f9",
  1498 => x"4f2648c0",
  1499 => x"78452080",
  1500 => x"80007469",
  1501 => x"63614220",
  1502 => x"10e9006b",
  1503 => x"2a990000",
  1504 => x"00000000",
  1505 => x"0010e900",
  1506 => x"002ab700",
  1507 => x"00000000",
  1508 => x"000010e9",
  1509 => x"00002ad5",
  1510 => x"e9000000",
  1511 => x"f3000010",
  1512 => x"0000002a",
  1513 => x"10e90000",
  1514 => x"2b110000",
  1515 => x"00000000",
  1516 => x"0010e900",
  1517 => x"002b2f00",
  1518 => x"00000000",
  1519 => x"000010e9",
  1520 => x"00002b4d",
  1521 => x"e9000000",
  1522 => x"00000010",
  1523 => x"00000000",
  1524 => x"117e0000",
  1525 => x"00000000",
  1526 => x"00000000",
  1527 => x"0017e100",
  1528 => x"534d4100",
  1529 => x"44415254",
  1530 => x"4d4f5220",
  1531 => x"616f4c00",
  1532 => x"2e2a2064",
  1533 => x"f0fe1e00",
  1534 => x"cd78c048",
  1535 => x"26097909",
  1536 => x"fe1e1e4f",
  1537 => x"487ebff0",
  1538 => x"1e4f2626",
  1539 => x"c148f0fe",
  1540 => x"1e4f2678",
  1541 => x"c048f0fe",
  1542 => x"1e4f2678",
  1543 => x"52c04a71",
  1544 => x"0e4f2652",
  1545 => x"5d5c5b5e",
  1546 => x"7186f40e",
  1547 => x"7e6d974d",
  1548 => x"974ca5c1",
  1549 => x"a6c8486c",
  1550 => x"c4486e58",
  1551 => x"c505a866",
  1552 => x"c048ff87",
  1553 => x"caff87e6",
  1554 => x"49a5c287",
  1555 => x"714b6c97",
  1556 => x"6b974ba3",
  1557 => x"7e6c974b",
  1558 => x"80c1486e",
  1559 => x"c758a6c8",
  1560 => x"58a6cc98",
  1561 => x"fe7c9770",
  1562 => x"487387e1",
  1563 => x"4d268ef4",
  1564 => x"4b264c26",
  1565 => x"5e0e4f26",
  1566 => x"f40e5c5b",
  1567 => x"d84c7186",
  1568 => x"ffc34a66",
  1569 => x"4ba4c29a",
  1570 => x"73496c97",
  1571 => x"517249a1",
  1572 => x"6e7e6c97",
  1573 => x"c880c148",
  1574 => x"98c758a6",
  1575 => x"7058a6cc",
  1576 => x"ff8ef454",
  1577 => x"1e1e87ca",
  1578 => x"e087e8fd",
  1579 => x"c0494abf",
  1580 => x"0299c0e0",
  1581 => x"1e7287cb",
  1582 => x"49ebedc2",
  1583 => x"c487f7fe",
  1584 => x"87fdfc86",
  1585 => x"c2fd7e70",
  1586 => x"4f262687",
  1587 => x"ebedc21e",
  1588 => x"87c7fd49",
  1589 => x"49e6e2c1",
  1590 => x"c587dafc",
  1591 => x"4f2687d9",
  1592 => x"5c5b5e0e",
  1593 => x"eec20e5d",
  1594 => x"c14abfca",
  1595 => x"49bff4e4",
  1596 => x"71bc724c",
  1597 => x"87dbfc4d",
  1598 => x"49744bc0",
  1599 => x"d50299d0",
  1600 => x"d0497587",
  1601 => x"c01e7199",
  1602 => x"c6ebc11e",
  1603 => x"1282734a",
  1604 => x"87e4c049",
  1605 => x"2cc186c8",
  1606 => x"abc8832d",
  1607 => x"87daff04",
  1608 => x"c187e8fb",
  1609 => x"c248f4e4",
  1610 => x"78bfcaee",
  1611 => x"4c264d26",
  1612 => x"4f264b26",
  1613 => x"00000000",
  1614 => x"48d0ff1e",
  1615 => x"ff78e1c8",
  1616 => x"78c548d4",
  1617 => x"c30266c4",
  1618 => x"78e0c387",
  1619 => x"c60266c8",
  1620 => x"48d4ff87",
  1621 => x"ff78f0c3",
  1622 => x"787148d4",
  1623 => x"c848d0ff",
  1624 => x"e0c078e1",
  1625 => x"0e4f2678",
  1626 => x"0e5c5b5e",
  1627 => x"edc24c71",
  1628 => x"eefa49eb",
  1629 => x"c04a7087",
  1630 => x"c204aab7",
  1631 => x"e0c387e3",
  1632 => x"87c905aa",
  1633 => x"48eae8c1",
  1634 => x"d4c278c1",
  1635 => x"aaf0c387",
  1636 => x"c187c905",
  1637 => x"c148e6e8",
  1638 => x"87f5c178",
  1639 => x"bfeae8c1",
  1640 => x"7287c702",
  1641 => x"b3c0c24b",
  1642 => x"4b7287c2",
  1643 => x"d1059c74",
  1644 => x"e6e8c187",
  1645 => x"e8c11ebf",
  1646 => x"721ebfea",
  1647 => x"87f8fd49",
  1648 => x"e8c186c8",
  1649 => x"c002bfe6",
  1650 => x"497387e0",
  1651 => x"9129b7c4",
  1652 => x"81c6eac1",
  1653 => x"9acf4a73",
  1654 => x"48c192c2",
  1655 => x"4a703072",
  1656 => x"4872baff",
  1657 => x"79709869",
  1658 => x"497387db",
  1659 => x"9129b7c4",
  1660 => x"81c6eac1",
  1661 => x"9acf4a73",
  1662 => x"48c392c2",
  1663 => x"4a703072",
  1664 => x"70b06948",
  1665 => x"eae8c179",
  1666 => x"c178c048",
  1667 => x"c048e6e8",
  1668 => x"ebedc278",
  1669 => x"87cbf849",
  1670 => x"b7c04a70",
  1671 => x"ddfd03aa",
  1672 => x"fc48c087",
  1673 => x"000087c8",
  1674 => x"00000000",
  1675 => x"711e0000",
  1676 => x"f2fc494a",
  1677 => x"1e4f2687",
  1678 => x"49724ac0",
  1679 => x"eac191c4",
  1680 => x"79c081c6",
  1681 => x"b7d082c1",
  1682 => x"87ee04aa",
  1683 => x"5e0e4f26",
  1684 => x"0e5d5c5b",
  1685 => x"faf64d71",
  1686 => x"c44a7587",
  1687 => x"c1922ab7",
  1688 => x"7582c6ea",
  1689 => x"c29ccf4c",
  1690 => x"4b496a94",
  1691 => x"9bc32b74",
  1692 => x"307448c2",
  1693 => x"bcff4c70",
  1694 => x"98714874",
  1695 => x"caf67a70",
  1696 => x"fa487387",
  1697 => x"000087e6",
  1698 => x"00000000",
  1699 => x"00000000",
  1700 => x"00000000",
  1701 => x"00000000",
  1702 => x"00000000",
  1703 => x"00000000",
  1704 => x"00000000",
  1705 => x"00000000",
  1706 => x"00000000",
  1707 => x"00000000",
  1708 => x"00000000",
  1709 => x"00000000",
  1710 => x"00000000",
  1711 => x"00000000",
  1712 => x"00000000",
  1713 => x"1e160000",
  1714 => x"362e2526",
  1715 => x"ff1e3e3d",
  1716 => x"e1c848d0",
  1717 => x"ff487178",
  1718 => x"267808d4",
  1719 => x"d0ff1e4f",
  1720 => x"78e1c848",
  1721 => x"d4ff4871",
  1722 => x"66c47808",
  1723 => x"08d4ff48",
  1724 => x"1e4f2678",
  1725 => x"66c44a71",
  1726 => x"49721e49",
  1727 => x"ff87deff",
  1728 => x"e0c048d0",
  1729 => x"4f262678",
  1730 => x"c44a711e",
  1731 => x"e0c11e66",
  1732 => x"c8ff49a2",
  1733 => x"4966c887",
  1734 => x"ff29b7c8",
  1735 => x"787148d4",
  1736 => x"c048d0ff",
  1737 => x"262678e0",
  1738 => x"d4ff1e4f",
  1739 => x"7affc34a",
  1740 => x"c848d0ff",
  1741 => x"7ade78e1",
  1742 => x"bff5edc2",
  1743 => x"c848497a",
  1744 => x"717a7028",
  1745 => x"7028d048",
  1746 => x"d848717a",
  1747 => x"ff7a7028",
  1748 => x"e0c048d0",
  1749 => x"0e4f2678",
  1750 => x"5d5c5b5e",
  1751 => x"c24c710e",
  1752 => x"4dbff5ed",
  1753 => x"d02b744b",
  1754 => x"83c19b66",
  1755 => x"04ab66d4",
  1756 => x"4bc087c2",
  1757 => x"66d04a74",
  1758 => x"ff317249",
  1759 => x"739975b9",
  1760 => x"70307248",
  1761 => x"b071484a",
  1762 => x"58f9edc2",
  1763 => x"2687dafe",
  1764 => x"264c264d",
  1765 => x"1e4f264b",
  1766 => x"c848d0ff",
  1767 => x"487178c9",
  1768 => x"7808d4ff",
  1769 => x"711e4f26",
  1770 => x"87eb494a",
  1771 => x"c848d0ff",
  1772 => x"1e4f2678",
  1773 => x"4b711e73",
  1774 => x"bfc5eec2",
  1775 => x"c287c302",
  1776 => x"d0ff87eb",
  1777 => x"78c9c848",
  1778 => x"e0c04973",
  1779 => x"48d4ffb1",
  1780 => x"edc27871",
  1781 => x"78c048f9",
  1782 => x"c50266c8",
  1783 => x"49ffc387",
  1784 => x"49c087c2",
  1785 => x"59c1eec2",
  1786 => x"c60266cc",
  1787 => x"d5d5c587",
  1788 => x"cf87c44a",
  1789 => x"c24affff",
  1790 => x"c25ac5ee",
  1791 => x"c148c5ee",
  1792 => x"2687c478",
  1793 => x"264c264d",
  1794 => x"0e4f264b",
  1795 => x"5d5c5b5e",
  1796 => x"c24a710e",
  1797 => x"4cbfc1ee",
  1798 => x"cb029a72",
  1799 => x"91c84987",
  1800 => x"4be9eec1",
  1801 => x"87c48371",
  1802 => x"4be9f2c1",
  1803 => x"49134dc0",
  1804 => x"edc29974",
  1805 => x"ffb9bffd",
  1806 => x"787148d4",
  1807 => x"852cb7c1",
  1808 => x"04adb7c8",
  1809 => x"edc287e8",
  1810 => x"c848bff9",
  1811 => x"fdedc280",
  1812 => x"87effe58",
  1813 => x"711e731e",
  1814 => x"9a4a134b",
  1815 => x"7287cb02",
  1816 => x"87e7fe49",
  1817 => x"059a4a13",
  1818 => x"dafe87f5",
  1819 => x"edc21e87",
  1820 => x"c249bff9",
  1821 => x"c148f9ed",
  1822 => x"c0c478a1",
  1823 => x"db03a9b7",
  1824 => x"48d4ff87",
  1825 => x"bffdedc2",
  1826 => x"f9edc278",
  1827 => x"edc249bf",
  1828 => x"a1c148f9",
  1829 => x"b7c0c478",
  1830 => x"87e504a9",
  1831 => x"c848d0ff",
  1832 => x"c5eec278",
  1833 => x"2678c048",
  1834 => x"0000004f",
  1835 => x"00000000",
  1836 => x"00000000",
  1837 => x"00005f5f",
  1838 => x"03030000",
  1839 => x"00030300",
  1840 => x"7f7f1400",
  1841 => x"147f7f14",
  1842 => x"2e240000",
  1843 => x"123a6b6b",
  1844 => x"366a4c00",
  1845 => x"32566c18",
  1846 => x"4f7e3000",
  1847 => x"683a7759",
  1848 => x"04000040",
  1849 => x"00000307",
  1850 => x"1c000000",
  1851 => x"0041633e",
  1852 => x"41000000",
  1853 => x"001c3e63",
  1854 => x"3e2a0800",
  1855 => x"2a3e1c1c",
  1856 => x"08080008",
  1857 => x"08083e3e",
  1858 => x"80000000",
  1859 => x"000060e0",
  1860 => x"08080000",
  1861 => x"08080808",
  1862 => x"00000000",
  1863 => x"00006060",
  1864 => x"30604000",
  1865 => x"03060c18",
  1866 => x"7f3e0001",
  1867 => x"3e7f4d59",
  1868 => x"06040000",
  1869 => x"00007f7f",
  1870 => x"63420000",
  1871 => x"464f5971",
  1872 => x"63220000",
  1873 => x"367f4949",
  1874 => x"161c1800",
  1875 => x"107f7f13",
  1876 => x"67270000",
  1877 => x"397d4545",
  1878 => x"7e3c0000",
  1879 => x"3079494b",
  1880 => x"01010000",
  1881 => x"070f7971",
  1882 => x"7f360000",
  1883 => x"367f4949",
  1884 => x"4f060000",
  1885 => x"1e3f6949",
  1886 => x"00000000",
  1887 => x"00006666",
  1888 => x"80000000",
  1889 => x"000066e6",
  1890 => x"08080000",
  1891 => x"22221414",
  1892 => x"14140000",
  1893 => x"14141414",
  1894 => x"22220000",
  1895 => x"08081414",
  1896 => x"03020000",
  1897 => x"060f5951",
  1898 => x"417f3e00",
  1899 => x"1e1f555d",
  1900 => x"7f7e0000",
  1901 => x"7e7f0909",
  1902 => x"7f7f0000",
  1903 => x"367f4949",
  1904 => x"3e1c0000",
  1905 => x"41414163",
  1906 => x"7f7f0000",
  1907 => x"1c3e6341",
  1908 => x"7f7f0000",
  1909 => x"41414949",
  1910 => x"7f7f0000",
  1911 => x"01010909",
  1912 => x"7f3e0000",
  1913 => x"7a7b4941",
  1914 => x"7f7f0000",
  1915 => x"7f7f0808",
  1916 => x"41000000",
  1917 => x"00417f7f",
  1918 => x"60200000",
  1919 => x"3f7f4040",
  1920 => x"087f7f00",
  1921 => x"4163361c",
  1922 => x"7f7f0000",
  1923 => x"40404040",
  1924 => x"067f7f00",
  1925 => x"7f7f060c",
  1926 => x"067f7f00",
  1927 => x"7f7f180c",
  1928 => x"7f3e0000",
  1929 => x"3e7f4141",
  1930 => x"7f7f0000",
  1931 => x"060f0909",
  1932 => x"417f3e00",
  1933 => x"407e7f61",
  1934 => x"7f7f0000",
  1935 => x"667f1909",
  1936 => x"6f260000",
  1937 => x"327b594d",
  1938 => x"01010000",
  1939 => x"01017f7f",
  1940 => x"7f3f0000",
  1941 => x"3f7f4040",
  1942 => x"3f0f0000",
  1943 => x"0f3f7070",
  1944 => x"307f7f00",
  1945 => x"7f7f3018",
  1946 => x"36634100",
  1947 => x"63361c1c",
  1948 => x"06030141",
  1949 => x"03067c7c",
  1950 => x"59716101",
  1951 => x"4143474d",
  1952 => x"7f000000",
  1953 => x"0041417f",
  1954 => x"06030100",
  1955 => x"6030180c",
  1956 => x"41000040",
  1957 => x"007f7f41",
  1958 => x"060c0800",
  1959 => x"080c0603",
  1960 => x"80808000",
  1961 => x"80808080",
  1962 => x"00000000",
  1963 => x"00040703",
  1964 => x"74200000",
  1965 => x"787c5454",
  1966 => x"7f7f0000",
  1967 => x"387c4444",
  1968 => x"7c380000",
  1969 => x"00444444",
  1970 => x"7c380000",
  1971 => x"7f7f4444",
  1972 => x"7c380000",
  1973 => x"185c5454",
  1974 => x"7e040000",
  1975 => x"0005057f",
  1976 => x"bc180000",
  1977 => x"7cfca4a4",
  1978 => x"7f7f0000",
  1979 => x"787c0404",
  1980 => x"00000000",
  1981 => x"00407d3d",
  1982 => x"80800000",
  1983 => x"007dfd80",
  1984 => x"7f7f0000",
  1985 => x"446c3810",
  1986 => x"00000000",
  1987 => x"00407f3f",
  1988 => x"0c7c7c00",
  1989 => x"787c0c18",
  1990 => x"7c7c0000",
  1991 => x"787c0404",
  1992 => x"7c380000",
  1993 => x"387c4444",
  1994 => x"fcfc0000",
  1995 => x"183c2424",
  1996 => x"3c180000",
  1997 => x"fcfc2424",
  1998 => x"7c7c0000",
  1999 => x"080c0404",
  2000 => x"5c480000",
  2001 => x"20745454",
  2002 => x"3f040000",
  2003 => x"0044447f",
  2004 => x"7c3c0000",
  2005 => x"7c7c4040",
  2006 => x"3c1c0000",
  2007 => x"1c3c6060",
  2008 => x"607c3c00",
  2009 => x"3c7c6030",
  2010 => x"386c4400",
  2011 => x"446c3810",
  2012 => x"bc1c0000",
  2013 => x"1c3c60e0",
  2014 => x"64440000",
  2015 => x"444c5c74",
  2016 => x"08080000",
  2017 => x"4141773e",
  2018 => x"00000000",
  2019 => x"00007f7f",
  2020 => x"41410000",
  2021 => x"08083e77",
  2022 => x"01010200",
  2023 => x"01020203",
  2024 => x"7f7f7f00",
  2025 => x"7f7f7f7f",
  2026 => x"1c080800",
  2027 => x"7f3e3e1c",
  2028 => x"3e7f7f7f",
  2029 => x"081c1c3e",
  2030 => x"18100008",
  2031 => x"10187c7c",
  2032 => x"30100000",
  2033 => x"10307c7c",
  2034 => x"60301000",
  2035 => x"061e7860",
  2036 => x"3c664200",
  2037 => x"42663c18",
  2038 => x"6a387800",
  2039 => x"386cc6c2",
  2040 => x"00006000",
  2041 => x"60000060",
  2042 => x"5b5e0e00",
  2043 => x"1e0e5d5c",
  2044 => x"eec24c71",
  2045 => x"c04dbfd6",
  2046 => x"741ec04b",
  2047 => x"87c702ab",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
