library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"c048a6c4",
     1 => x"c487c578",
     2 => x"78c148a6",
     3 => x"731e66c4",
     4 => x"87dfee49",
     5 => x"e0c086c8",
     6 => x"87efef49",
     7 => x"6a4aa5c4",
     8 => x"87f0f049",
     9 => x"cb87c6f1",
    10 => x"c883c185",
    11 => x"ff04abb7",
    12 => x"262687c7",
    13 => x"264c264d",
    14 => x"1e4f264b",
    15 => x"eec24a71",
    16 => x"eec25ada",
    17 => x"78c748da",
    18 => x"87ddfe49",
    19 => x"731e4f26",
    20 => x"c04a711e",
    21 => x"d303aab7",
    22 => x"dfcec287",
    23 => x"87c405bf",
    24 => x"87c24bc1",
    25 => x"cec24bc0",
    26 => x"87c45be3",
    27 => x"5ae3cec2",
    28 => x"bfdfcec2",
    29 => x"c19ac14a",
    30 => x"ec49a2c0",
    31 => x"48fc87e8",
    32 => x"bfdfcec2",
    33 => x"87effe78",
    34 => x"c44a711e",
    35 => x"49721e66",
    36 => x"2687f5e9",
    37 => x"c21e4f26",
    38 => x"49bfdfce",
    39 => x"c287cfe6",
    40 => x"e848ceee",
    41 => x"eec278bf",
    42 => x"bfec48ca",
    43 => x"ceeec278",
    44 => x"c3494abf",
    45 => x"b7c899ff",
    46 => x"7148722a",
    47 => x"d6eec2b0",
    48 => x"0e4f2658",
    49 => x"5d5c5b5e",
    50 => x"ff4b710e",
    51 => x"eec287c8",
    52 => x"50c048c9",
    53 => x"f5e54973",
    54 => x"4c497087",
    55 => x"eecb9cc2",
    56 => x"87c3cb49",
    57 => x"c24d4970",
    58 => x"bf97c9ee",
    59 => x"87e2c105",
    60 => x"c24966d0",
    61 => x"99bfd2ee",
    62 => x"d487d605",
    63 => x"eec24966",
    64 => x"0599bfca",
    65 => x"497387cb",
    66 => x"7087c3e5",
    67 => x"c1c10298",
    68 => x"fe4cc187",
    69 => x"497587c0",
    70 => x"7087d8ca",
    71 => x"87c60298",
    72 => x"48c9eec2",
    73 => x"eec250c1",
    74 => x"05bf97c9",
    75 => x"c287e3c0",
    76 => x"49bfd2ee",
    77 => x"059966d0",
    78 => x"c287d6ff",
    79 => x"49bfcaee",
    80 => x"059966d4",
    81 => x"7387caff",
    82 => x"87c2e449",
    83 => x"fe059870",
    84 => x"487487ff",
    85 => x"0e87dcfb",
    86 => x"5d5c5b5e",
    87 => x"c086f40e",
    88 => x"bfec4c4d",
    89 => x"48a6c47e",
    90 => x"bfd6eec2",
    91 => x"c01ec178",
    92 => x"fd49c71e",
    93 => x"86c887cd",
    94 => x"cd029870",
    95 => x"fb49ff87",
    96 => x"dac187cc",
    97 => x"87c6e349",
    98 => x"eec24dc1",
    99 => x"02bf97c9",
   100 => x"fed487c3",
   101 => x"ceeec287",
   102 => x"cec24bbf",
   103 => x"c005bfdf",
   104 => x"fdc387e9",
   105 => x"87e6e249",
   106 => x"e249fac3",
   107 => x"497387e0",
   108 => x"7199ffc3",
   109 => x"fb49c01e",
   110 => x"497387ce",
   111 => x"7129b7c8",
   112 => x"fb49c11e",
   113 => x"86c887c2",
   114 => x"c287fac5",
   115 => x"4bbfd2ee",
   116 => x"87dd029b",
   117 => x"bfdbcec2",
   118 => x"87d7c749",
   119 => x"c4059870",
   120 => x"d24bc087",
   121 => x"49e0c287",
   122 => x"c287fcc6",
   123 => x"c658dfce",
   124 => x"dbcec287",
   125 => x"7378c048",
   126 => x"0599c249",
   127 => x"ebc387cd",
   128 => x"87cae149",
   129 => x"99c24970",
   130 => x"fb87c202",
   131 => x"c149734c",
   132 => x"87cd0599",
   133 => x"e049f4c3",
   134 => x"497087f4",
   135 => x"c20299c2",
   136 => x"734cfa87",
   137 => x"0599c849",
   138 => x"f5c387cd",
   139 => x"87dee049",
   140 => x"99c24970",
   141 => x"c287d402",
   142 => x"02bfdaee",
   143 => x"c14887c9",
   144 => x"deeec288",
   145 => x"ff87c258",
   146 => x"734dc14c",
   147 => x"0599c449",
   148 => x"f2c387ce",
   149 => x"f5dfff49",
   150 => x"c2497087",
   151 => x"87db0299",
   152 => x"bfdaeec2",
   153 => x"b7c7487e",
   154 => x"87cb03a8",
   155 => x"80c1486e",
   156 => x"58deeec2",
   157 => x"fe87c2c0",
   158 => x"c34dc14c",
   159 => x"dfff49fd",
   160 => x"497087cc",
   161 => x"d50299c2",
   162 => x"daeec287",
   163 => x"c9c002bf",
   164 => x"daeec287",
   165 => x"c078c048",
   166 => x"4cfd87c2",
   167 => x"fac34dc1",
   168 => x"e9deff49",
   169 => x"c2497087",
   170 => x"87d90299",
   171 => x"bfdaeec2",
   172 => x"a8b7c748",
   173 => x"87c9c003",
   174 => x"48daeec2",
   175 => x"c2c078c7",
   176 => x"c14cfc87",
   177 => x"acb7c04d",
   178 => x"87d1c003",
   179 => x"c14a66c4",
   180 => x"026a82d8",
   181 => x"6a87c6c0",
   182 => x"7349744b",
   183 => x"c31ec00f",
   184 => x"dac11ef0",
   185 => x"87dbf749",
   186 => x"987086c8",
   187 => x"87e2c002",
   188 => x"c248a6c8",
   189 => x"78bfdaee",
   190 => x"cb4966c8",
   191 => x"4866c491",
   192 => x"7e708071",
   193 => x"c002bf6e",
   194 => x"bf6e87c8",
   195 => x"4966c84b",
   196 => x"9d750f73",
   197 => x"87c8c002",
   198 => x"bfdaeec2",
   199 => x"87c9f349",
   200 => x"bfe3cec2",
   201 => x"87ddc002",
   202 => x"87c7c249",
   203 => x"c0029870",
   204 => x"eec287d3",
   205 => x"f249bfda",
   206 => x"49c087ef",
   207 => x"c287cff4",
   208 => x"c048e3ce",
   209 => x"f38ef478",
   210 => x"5e0e87e9",
   211 => x"0e5d5c5b",
   212 => x"c24c711e",
   213 => x"49bfd6ee",
   214 => x"4da1cdc1",
   215 => x"6981d1c1",
   216 => x"029c747e",
   217 => x"a5c487cf",
   218 => x"c27b744b",
   219 => x"49bfd6ee",
   220 => x"6e87c8f3",
   221 => x"059c747b",
   222 => x"4bc087c4",
   223 => x"4bc187c2",
   224 => x"c9f34973",
   225 => x"0266d487",
   226 => x"da4987c7",
   227 => x"c24a7087",
   228 => x"c24ac087",
   229 => x"265ae7ce",
   230 => x"0087d8f2",
   231 => x"00000000",
   232 => x"00000000",
   233 => x"1e000000",
   234 => x"c8ff4a71",
   235 => x"a17249bf",
   236 => x"1e4f2648",
   237 => x"89bfc8ff",
   238 => x"c0c0c0fe",
   239 => x"01a9c0c0",
   240 => x"4ac087c4",
   241 => x"4ac187c2",
   242 => x"4f264872",
   243 => x"5c5b5e0e",
   244 => x"4b710e5d",
   245 => x"d04cd4ff",
   246 => x"78c04866",
   247 => x"dbff49d6",
   248 => x"ffc387ec",
   249 => x"c3496c7c",
   250 => x"4d7199ff",
   251 => x"99f0c349",
   252 => x"05a9e0c1",
   253 => x"ffc387cb",
   254 => x"c3486c7c",
   255 => x"0866d098",
   256 => x"7cffc378",
   257 => x"c8494a6c",
   258 => x"7cffc331",
   259 => x"b2714a6c",
   260 => x"31c84972",
   261 => x"6c7cffc3",
   262 => x"72b2714a",
   263 => x"c331c849",
   264 => x"4a6c7cff",
   265 => x"d0ffb271",
   266 => x"78e0c048",
   267 => x"c2029b73",
   268 => x"757b7287",
   269 => x"264d2648",
   270 => x"264b264c",
   271 => x"4f261e4f",
   272 => x"5c5b5e0e",
   273 => x"7686f80e",
   274 => x"49a6c81e",
   275 => x"c487fdfd",
   276 => x"6e4b7086",
   277 => x"03a8c248",
   278 => x"7387c6c3",
   279 => x"9af0c34a",
   280 => x"02aad0c1",
   281 => x"e0c187c7",
   282 => x"f4c205aa",
   283 => x"c8497387",
   284 => x"87c30299",
   285 => x"7387c6ff",
   286 => x"c29cc34c",
   287 => x"cdc105ac",
   288 => x"4966c487",
   289 => x"1e7131c9",
   290 => x"d44a66c4",
   291 => x"deeec292",
   292 => x"fe817249",
   293 => x"c487d8d4",
   294 => x"c01e4966",
   295 => x"d9ff49e3",
   296 => x"49d887d1",
   297 => x"87e6d8ff",
   298 => x"c21ec0c8",
   299 => x"fd49cedd",
   300 => x"ff87e8f0",
   301 => x"e0c048d0",
   302 => x"ceddc278",
   303 => x"4a66d01e",
   304 => x"eec292d4",
   305 => x"817249de",
   306 => x"87e0d2fe",
   307 => x"acc186d0",
   308 => x"87cdc105",
   309 => x"c94966c4",
   310 => x"c41e7131",
   311 => x"92d44a66",
   312 => x"49deeec2",
   313 => x"d3fe8172",
   314 => x"ddc287c5",
   315 => x"66c81ece",
   316 => x"c292d44a",
   317 => x"7249deee",
   318 => x"ecd0fe81",
   319 => x"4966c887",
   320 => x"49e3c01e",
   321 => x"87ebd7ff",
   322 => x"d7ff49d7",
   323 => x"c0c887c0",
   324 => x"ceddc21e",
   325 => x"eceefd49",
   326 => x"ff86d087",
   327 => x"e0c048d0",
   328 => x"fc8ef878",
   329 => x"5e0e87d1",
   330 => x"0e5d5c5b",
   331 => x"ff4d711e",
   332 => x"66d44cd4",
   333 => x"b7c3487e",
   334 => x"87c506a8",
   335 => x"e2c148c0",
   336 => x"fe497587",
   337 => x"7587f9e0",
   338 => x"4b66c41e",
   339 => x"eec293d4",
   340 => x"497383de",
   341 => x"87f5cbfe",
   342 => x"4b6b83c8",
   343 => x"c848d0ff",
   344 => x"7cdd78e1",
   345 => x"ffc34973",
   346 => x"737c7199",
   347 => x"29b7c849",
   348 => x"7199ffc3",
   349 => x"d049737c",
   350 => x"ffc329b7",
   351 => x"737c7199",
   352 => x"29b7d849",
   353 => x"7cc07c71",
   354 => x"7c7c7c7c",
   355 => x"7c7c7c7c",
   356 => x"c07c7c7c",
   357 => x"66c478e0",
   358 => x"ff49dc1e",
   359 => x"c887d4d5",
   360 => x"26487386",
   361 => x"0e87cefa",
   362 => x"5d5c5b5e",
   363 => x"7e711e0e",
   364 => x"6e4bd4ff",
   365 => x"c6efc21e",
   366 => x"d0cafe49",
   367 => x"7086c487",
   368 => x"c3029d4d",
   369 => x"efc287c3",
   370 => x"6e4cbfce",
   371 => x"efdefe49",
   372 => x"48d0ff87",
   373 => x"c178c5c8",
   374 => x"4ac07bd6",
   375 => x"82c17b15",
   376 => x"aab7e0c0",
   377 => x"ff87f504",
   378 => x"78c448d0",
   379 => x"c178c5c8",
   380 => x"7bc17bd3",
   381 => x"9c7478c4",
   382 => x"87fcc102",
   383 => x"7eceddc2",
   384 => x"8c4dc0c8",
   385 => x"03acb7c0",
   386 => x"c0c887c6",
   387 => x"4cc04da4",
   388 => x"97ffe9c2",
   389 => x"99d049bf",
   390 => x"c087d202",
   391 => x"c6efc21e",
   392 => x"c4ccfe49",
   393 => x"7086c487",
   394 => x"efc04a49",
   395 => x"ceddc287",
   396 => x"c6efc21e",
   397 => x"f0cbfe49",
   398 => x"7086c487",
   399 => x"d0ff4a49",
   400 => x"78c5c848",
   401 => x"6e7bd4c1",
   402 => x"6e7bbf97",
   403 => x"7080c148",
   404 => x"058dc17e",
   405 => x"ff87f0ff",
   406 => x"78c448d0",
   407 => x"c5059a72",
   408 => x"c048c087",
   409 => x"1ec187e5",
   410 => x"49c6efc2",
   411 => x"87d8c9fe",
   412 => x"9c7486c4",
   413 => x"87c4fe05",
   414 => x"c848d0ff",
   415 => x"d3c178c5",
   416 => x"c47bc07b",
   417 => x"c248c178",
   418 => x"2648c087",
   419 => x"4c264d26",
   420 => x"4f264b26",
   421 => x"5c5b5e0e",
   422 => x"cc4b710e",
   423 => x"87d80266",
   424 => x"8cf0c04c",
   425 => x"7487d802",
   426 => x"028ac14a",
   427 => x"028a87d1",
   428 => x"028a87cd",
   429 => x"87d787c9",
   430 => x"eafb4973",
   431 => x"7487d087",
   432 => x"f949c01e",
   433 => x"1e7487e0",
   434 => x"d9f94973",
   435 => x"fe86c887",
   436 => x"1e0087fc",
   437 => x"bfe1dcc2",
   438 => x"c2b9c149",
   439 => x"ff59e5dc",
   440 => x"ffc348d4",
   441 => x"48d0ff78",
   442 => x"ff78e1c8",
   443 => x"78c148d4",
   444 => x"787131c4",
   445 => x"c048d0ff",
   446 => x"4f2678e0",
   447 => x"d5dcc21e",
   448 => x"c6efc21e",
   449 => x"c4c5fe49",
   450 => x"7086c487",
   451 => x"87c30298",
   452 => x"2687c0ff",
   453 => x"4b35314f",
   454 => x"20205a48",
   455 => x"47464320",
   456 => x"00000000",
   457 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
