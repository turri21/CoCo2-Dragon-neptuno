
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"dc",x"ef",x"c2",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"dc",x"ef",x"c2"),
    14 => (x"48",x"e8",x"dc",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"cb",x"dc"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"48",x"11",x"1e",x"4f"),
    50 => (x"78",x"08",x"d4",x"ff"),
    51 => (x"c1",x"48",x"66",x"c4"),
    52 => (x"58",x"a6",x"c8",x"88"),
    53 => (x"ed",x"05",x"98",x"70"),
    54 => (x"1e",x"4f",x"26",x"87"),
    55 => (x"c3",x"48",x"d4",x"ff"),
    56 => (x"51",x"68",x"78",x"ff"),
    57 => (x"c1",x"48",x"66",x"c4"),
    58 => (x"58",x"a6",x"c8",x"88"),
    59 => (x"eb",x"05",x"98",x"70"),
    60 => (x"1e",x"4f",x"26",x"87"),
    61 => (x"d4",x"ff",x"1e",x"73"),
    62 => (x"7b",x"ff",x"c3",x"4b"),
    63 => (x"ff",x"c3",x"4a",x"6b"),
    64 => (x"c8",x"49",x"6b",x"7b"),
    65 => (x"c3",x"b1",x"72",x"32"),
    66 => (x"4a",x"6b",x"7b",x"ff"),
    67 => (x"b2",x"71",x"31",x"c8"),
    68 => (x"6b",x"7b",x"ff",x"c3"),
    69 => (x"72",x"32",x"c8",x"49"),
    70 => (x"c4",x"48",x"71",x"b1"),
    71 => (x"26",x"4d",x"26",x"87"),
    72 => (x"26",x"4b",x"26",x"4c"),
    73 => (x"5b",x"5e",x"0e",x"4f"),
    74 => (x"71",x"0e",x"5d",x"5c"),
    75 => (x"4c",x"d4",x"ff",x"4a"),
    76 => (x"ff",x"c3",x"49",x"72"),
    77 => (x"c2",x"7c",x"71",x"99"),
    78 => (x"05",x"bf",x"e8",x"dc"),
    79 => (x"66",x"d0",x"87",x"c8"),
    80 => (x"d4",x"30",x"c9",x"48"),
    81 => (x"66",x"d0",x"58",x"a6"),
    82 => (x"c3",x"29",x"d8",x"49"),
    83 => (x"7c",x"71",x"99",x"ff"),
    84 => (x"d0",x"49",x"66",x"d0"),
    85 => (x"99",x"ff",x"c3",x"29"),
    86 => (x"66",x"d0",x"7c",x"71"),
    87 => (x"c3",x"29",x"c8",x"49"),
    88 => (x"7c",x"71",x"99",x"ff"),
    89 => (x"c3",x"49",x"66",x"d0"),
    90 => (x"7c",x"71",x"99",x"ff"),
    91 => (x"29",x"d0",x"49",x"72"),
    92 => (x"71",x"99",x"ff",x"c3"),
    93 => (x"c9",x"4b",x"6c",x"7c"),
    94 => (x"c3",x"4d",x"ff",x"f0"),
    95 => (x"d0",x"05",x"ab",x"ff"),
    96 => (x"7c",x"ff",x"c3",x"87"),
    97 => (x"8d",x"c1",x"4b",x"6c"),
    98 => (x"c3",x"87",x"c6",x"02"),
    99 => (x"f0",x"02",x"ab",x"ff"),
   100 => (x"fe",x"48",x"73",x"87"),
   101 => (x"c0",x"1e",x"87",x"c7"),
   102 => (x"48",x"d4",x"ff",x"49"),
   103 => (x"c1",x"78",x"ff",x"c3"),
   104 => (x"b7",x"c8",x"c3",x"81"),
   105 => (x"87",x"f1",x"04",x"a9"),
   106 => (x"73",x"1e",x"4f",x"26"),
   107 => (x"c4",x"87",x"e7",x"1e"),
   108 => (x"c0",x"4b",x"df",x"f8"),
   109 => (x"f0",x"ff",x"c0",x"1e"),
   110 => (x"fd",x"49",x"f7",x"c1"),
   111 => (x"86",x"c4",x"87",x"e7"),
   112 => (x"c0",x"05",x"a8",x"c1"),
   113 => (x"d4",x"ff",x"87",x"ea"),
   114 => (x"78",x"ff",x"c3",x"48"),
   115 => (x"c0",x"c0",x"c0",x"c1"),
   116 => (x"c0",x"1e",x"c0",x"c0"),
   117 => (x"e9",x"c1",x"f0",x"e1"),
   118 => (x"87",x"c9",x"fd",x"49"),
   119 => (x"98",x"70",x"86",x"c4"),
   120 => (x"ff",x"87",x"ca",x"05"),
   121 => (x"ff",x"c3",x"48",x"d4"),
   122 => (x"cb",x"48",x"c1",x"78"),
   123 => (x"87",x"e6",x"fe",x"87"),
   124 => (x"fe",x"05",x"8b",x"c1"),
   125 => (x"48",x"c0",x"87",x"fd"),
   126 => (x"1e",x"87",x"e6",x"fc"),
   127 => (x"d4",x"ff",x"1e",x"73"),
   128 => (x"78",x"ff",x"c3",x"48"),
   129 => (x"1e",x"c0",x"4b",x"d3"),
   130 => (x"c1",x"f0",x"ff",x"c0"),
   131 => (x"d4",x"fc",x"49",x"c1"),
   132 => (x"70",x"86",x"c4",x"87"),
   133 => (x"87",x"ca",x"05",x"98"),
   134 => (x"c3",x"48",x"d4",x"ff"),
   135 => (x"48",x"c1",x"78",x"ff"),
   136 => (x"f1",x"fd",x"87",x"cb"),
   137 => (x"05",x"8b",x"c1",x"87"),
   138 => (x"c0",x"87",x"db",x"ff"),
   139 => (x"87",x"f1",x"fb",x"48"),
   140 => (x"5c",x"5b",x"5e",x"0e"),
   141 => (x"4c",x"d4",x"ff",x"0e"),
   142 => (x"c6",x"87",x"db",x"fd"),
   143 => (x"e1",x"c0",x"1e",x"ea"),
   144 => (x"49",x"c8",x"c1",x"f0"),
   145 => (x"c4",x"87",x"de",x"fb"),
   146 => (x"02",x"a8",x"c1",x"86"),
   147 => (x"ea",x"fe",x"87",x"c8"),
   148 => (x"c1",x"48",x"c0",x"87"),
   149 => (x"da",x"fa",x"87",x"e2"),
   150 => (x"cf",x"49",x"70",x"87"),
   151 => (x"c6",x"99",x"ff",x"ff"),
   152 => (x"c8",x"02",x"a9",x"ea"),
   153 => (x"87",x"d3",x"fe",x"87"),
   154 => (x"cb",x"c1",x"48",x"c0"),
   155 => (x"7c",x"ff",x"c3",x"87"),
   156 => (x"fc",x"4b",x"f1",x"c0"),
   157 => (x"98",x"70",x"87",x"f4"),
   158 => (x"87",x"eb",x"c0",x"02"),
   159 => (x"ff",x"c0",x"1e",x"c0"),
   160 => (x"49",x"fa",x"c1",x"f0"),
   161 => (x"c4",x"87",x"de",x"fa"),
   162 => (x"05",x"98",x"70",x"86"),
   163 => (x"ff",x"c3",x"87",x"d9"),
   164 => (x"c3",x"49",x"6c",x"7c"),
   165 => (x"7c",x"7c",x"7c",x"ff"),
   166 => (x"99",x"c0",x"c1",x"7c"),
   167 => (x"c1",x"87",x"c4",x"02"),
   168 => (x"c0",x"87",x"d5",x"48"),
   169 => (x"c2",x"87",x"d1",x"48"),
   170 => (x"87",x"c4",x"05",x"ab"),
   171 => (x"87",x"c8",x"48",x"c0"),
   172 => (x"fe",x"05",x"8b",x"c1"),
   173 => (x"48",x"c0",x"87",x"fd"),
   174 => (x"1e",x"87",x"e4",x"f9"),
   175 => (x"dc",x"c2",x"1e",x"73"),
   176 => (x"78",x"c1",x"48",x"e8"),
   177 => (x"d0",x"ff",x"4b",x"c7"),
   178 => (x"fb",x"78",x"c2",x"48"),
   179 => (x"d0",x"ff",x"87",x"c8"),
   180 => (x"c0",x"78",x"c3",x"48"),
   181 => (x"d0",x"e5",x"c0",x"1e"),
   182 => (x"f9",x"49",x"c0",x"c1"),
   183 => (x"86",x"c4",x"87",x"c7"),
   184 => (x"c1",x"05",x"a8",x"c1"),
   185 => (x"ab",x"c2",x"4b",x"87"),
   186 => (x"c0",x"87",x"c5",x"05"),
   187 => (x"87",x"f9",x"c0",x"48"),
   188 => (x"ff",x"05",x"8b",x"c1"),
   189 => (x"f7",x"fc",x"87",x"d0"),
   190 => (x"ec",x"dc",x"c2",x"87"),
   191 => (x"05",x"98",x"70",x"58"),
   192 => (x"1e",x"c1",x"87",x"cd"),
   193 => (x"c1",x"f0",x"ff",x"c0"),
   194 => (x"d8",x"f8",x"49",x"d0"),
   195 => (x"ff",x"86",x"c4",x"87"),
   196 => (x"ff",x"c3",x"48",x"d4"),
   197 => (x"87",x"e0",x"c4",x"78"),
   198 => (x"58",x"f0",x"dc",x"c2"),
   199 => (x"c2",x"48",x"d0",x"ff"),
   200 => (x"48",x"d4",x"ff",x"78"),
   201 => (x"c1",x"78",x"ff",x"c3"),
   202 => (x"87",x"f5",x"f7",x"48"),
   203 => (x"5c",x"5b",x"5e",x"0e"),
   204 => (x"4a",x"71",x"0e",x"5d"),
   205 => (x"ff",x"4d",x"ff",x"c3"),
   206 => (x"7c",x"75",x"4c",x"d4"),
   207 => (x"c4",x"48",x"d0",x"ff"),
   208 => (x"7c",x"75",x"78",x"c3"),
   209 => (x"ff",x"c0",x"1e",x"72"),
   210 => (x"49",x"d8",x"c1",x"f0"),
   211 => (x"c4",x"87",x"d6",x"f7"),
   212 => (x"02",x"98",x"70",x"86"),
   213 => (x"48",x"c0",x"87",x"c5"),
   214 => (x"75",x"87",x"f0",x"c0"),
   215 => (x"7c",x"fe",x"c3",x"7c"),
   216 => (x"d4",x"1e",x"c0",x"c8"),
   217 => (x"dc",x"f5",x"49",x"66"),
   218 => (x"75",x"86",x"c4",x"87"),
   219 => (x"75",x"7c",x"75",x"7c"),
   220 => (x"e0",x"da",x"d8",x"7c"),
   221 => (x"6c",x"7c",x"75",x"4b"),
   222 => (x"c5",x"05",x"99",x"49"),
   223 => (x"05",x"8b",x"c1",x"87"),
   224 => (x"7c",x"75",x"87",x"f3"),
   225 => (x"c2",x"48",x"d0",x"ff"),
   226 => (x"f6",x"48",x"c1",x"78"),
   227 => (x"ff",x"1e",x"87",x"cf"),
   228 => (x"d0",x"ff",x"4a",x"d4"),
   229 => (x"78",x"d1",x"c4",x"48"),
   230 => (x"c1",x"7a",x"ff",x"c3"),
   231 => (x"87",x"f8",x"05",x"89"),
   232 => (x"73",x"1e",x"4f",x"26"),
   233 => (x"c5",x"4b",x"71",x"1e"),
   234 => (x"4a",x"df",x"cd",x"ee"),
   235 => (x"c3",x"48",x"d4",x"ff"),
   236 => (x"48",x"68",x"78",x"ff"),
   237 => (x"02",x"a8",x"fe",x"c3"),
   238 => (x"8a",x"c1",x"87",x"c5"),
   239 => (x"72",x"87",x"ed",x"05"),
   240 => (x"87",x"c5",x"05",x"9a"),
   241 => (x"ea",x"c0",x"48",x"c0"),
   242 => (x"02",x"9b",x"73",x"87"),
   243 => (x"66",x"c8",x"87",x"cc"),
   244 => (x"f4",x"49",x"73",x"1e"),
   245 => (x"86",x"c4",x"87",x"c5"),
   246 => (x"66",x"c8",x"87",x"c6"),
   247 => (x"87",x"ee",x"fe",x"49"),
   248 => (x"c3",x"48",x"d4",x"ff"),
   249 => (x"73",x"78",x"78",x"ff"),
   250 => (x"87",x"c5",x"05",x"9b"),
   251 => (x"d0",x"48",x"d0",x"ff"),
   252 => (x"f4",x"48",x"c1",x"78"),
   253 => (x"73",x"1e",x"87",x"eb"),
   254 => (x"c0",x"4a",x"71",x"1e"),
   255 => (x"48",x"d4",x"ff",x"4b"),
   256 => (x"ff",x"78",x"ff",x"c3"),
   257 => (x"c3",x"c4",x"48",x"d0"),
   258 => (x"48",x"d4",x"ff",x"78"),
   259 => (x"72",x"78",x"ff",x"c3"),
   260 => (x"f0",x"ff",x"c0",x"1e"),
   261 => (x"f4",x"49",x"d1",x"c1"),
   262 => (x"86",x"c4",x"87",x"cb"),
   263 => (x"cd",x"05",x"98",x"70"),
   264 => (x"1e",x"c0",x"c8",x"87"),
   265 => (x"fd",x"49",x"66",x"cc"),
   266 => (x"86",x"c4",x"87",x"f8"),
   267 => (x"d0",x"ff",x"4b",x"70"),
   268 => (x"73",x"78",x"c2",x"48"),
   269 => (x"87",x"e9",x"f3",x"48"),
   270 => (x"5c",x"5b",x"5e",x"0e"),
   271 => (x"1e",x"c0",x"0e",x"5d"),
   272 => (x"c1",x"f0",x"ff",x"c0"),
   273 => (x"dc",x"f3",x"49",x"c9"),
   274 => (x"c2",x"1e",x"d2",x"87"),
   275 => (x"fd",x"49",x"f0",x"dc"),
   276 => (x"86",x"c8",x"87",x"d0"),
   277 => (x"84",x"c1",x"4c",x"c0"),
   278 => (x"04",x"ac",x"b7",x"d2"),
   279 => (x"dc",x"c2",x"87",x"f8"),
   280 => (x"49",x"bf",x"97",x"f0"),
   281 => (x"c1",x"99",x"c0",x"c3"),
   282 => (x"c0",x"05",x"a9",x"c0"),
   283 => (x"dc",x"c2",x"87",x"e7"),
   284 => (x"49",x"bf",x"97",x"f7"),
   285 => (x"dc",x"c2",x"31",x"d0"),
   286 => (x"4a",x"bf",x"97",x"f8"),
   287 => (x"b1",x"72",x"32",x"c8"),
   288 => (x"97",x"f9",x"dc",x"c2"),
   289 => (x"71",x"b1",x"4a",x"bf"),
   290 => (x"ff",x"ff",x"cf",x"4c"),
   291 => (x"84",x"c1",x"9c",x"ff"),
   292 => (x"e7",x"c1",x"34",x"ca"),
   293 => (x"f9",x"dc",x"c2",x"87"),
   294 => (x"c1",x"49",x"bf",x"97"),
   295 => (x"c2",x"99",x"c6",x"31"),
   296 => (x"bf",x"97",x"fa",x"dc"),
   297 => (x"2a",x"b7",x"c7",x"4a"),
   298 => (x"dc",x"c2",x"b1",x"72"),
   299 => (x"4a",x"bf",x"97",x"f5"),
   300 => (x"c2",x"9d",x"cf",x"4d"),
   301 => (x"bf",x"97",x"f6",x"dc"),
   302 => (x"ca",x"9a",x"c3",x"4a"),
   303 => (x"f7",x"dc",x"c2",x"32"),
   304 => (x"c2",x"4b",x"bf",x"97"),
   305 => (x"c2",x"b2",x"73",x"33"),
   306 => (x"bf",x"97",x"f8",x"dc"),
   307 => (x"9b",x"c0",x"c3",x"4b"),
   308 => (x"73",x"2b",x"b7",x"c6"),
   309 => (x"c1",x"81",x"c2",x"b2"),
   310 => (x"70",x"30",x"71",x"48"),
   311 => (x"75",x"48",x"c1",x"49"),
   312 => (x"72",x"4d",x"70",x"30"),
   313 => (x"71",x"84",x"c1",x"4c"),
   314 => (x"b7",x"c0",x"c8",x"94"),
   315 => (x"87",x"cc",x"06",x"ad"),
   316 => (x"2d",x"b7",x"34",x"c1"),
   317 => (x"ad",x"b7",x"c0",x"c8"),
   318 => (x"87",x"f4",x"ff",x"01"),
   319 => (x"dc",x"f0",x"48",x"74"),
   320 => (x"5b",x"5e",x"0e",x"87"),
   321 => (x"f8",x"0e",x"5d",x"5c"),
   322 => (x"d6",x"e5",x"c2",x"86"),
   323 => (x"c2",x"78",x"c0",x"48"),
   324 => (x"c0",x"1e",x"ce",x"dd"),
   325 => (x"87",x"de",x"fb",x"49"),
   326 => (x"98",x"70",x"86",x"c4"),
   327 => (x"c0",x"87",x"c5",x"05"),
   328 => (x"87",x"ce",x"c9",x"48"),
   329 => (x"7e",x"c1",x"4d",x"c0"),
   330 => (x"bf",x"cb",x"f2",x"c0"),
   331 => (x"c4",x"de",x"c2",x"49"),
   332 => (x"4b",x"c8",x"71",x"4a"),
   333 => (x"70",x"87",x"f3",x"ec"),
   334 => (x"87",x"c2",x"05",x"98"),
   335 => (x"f2",x"c0",x"7e",x"c0"),
   336 => (x"c2",x"49",x"bf",x"c7"),
   337 => (x"71",x"4a",x"e0",x"de"),
   338 => (x"dd",x"ec",x"4b",x"c8"),
   339 => (x"05",x"98",x"70",x"87"),
   340 => (x"7e",x"c0",x"87",x"c2"),
   341 => (x"fd",x"c0",x"02",x"6e"),
   342 => (x"d4",x"e4",x"c2",x"87"),
   343 => (x"e5",x"c2",x"4d",x"bf"),
   344 => (x"7e",x"bf",x"9f",x"cc"),
   345 => (x"ea",x"d6",x"c5",x"48"),
   346 => (x"87",x"c7",x"05",x"a8"),
   347 => (x"bf",x"d4",x"e4",x"c2"),
   348 => (x"6e",x"87",x"ce",x"4d"),
   349 => (x"d5",x"e9",x"ca",x"48"),
   350 => (x"87",x"c5",x"02",x"a8"),
   351 => (x"f1",x"c7",x"48",x"c0"),
   352 => (x"ce",x"dd",x"c2",x"87"),
   353 => (x"f9",x"49",x"75",x"1e"),
   354 => (x"86",x"c4",x"87",x"ec"),
   355 => (x"c5",x"05",x"98",x"70"),
   356 => (x"c7",x"48",x"c0",x"87"),
   357 => (x"f2",x"c0",x"87",x"dc"),
   358 => (x"c2",x"49",x"bf",x"c7"),
   359 => (x"71",x"4a",x"e0",x"de"),
   360 => (x"c5",x"eb",x"4b",x"c8"),
   361 => (x"05",x"98",x"70",x"87"),
   362 => (x"e5",x"c2",x"87",x"c8"),
   363 => (x"78",x"c1",x"48",x"d6"),
   364 => (x"f2",x"c0",x"87",x"da"),
   365 => (x"c2",x"49",x"bf",x"cb"),
   366 => (x"71",x"4a",x"c4",x"de"),
   367 => (x"e9",x"ea",x"4b",x"c8"),
   368 => (x"02",x"98",x"70",x"87"),
   369 => (x"c0",x"87",x"c5",x"c0"),
   370 => (x"87",x"e6",x"c6",x"48"),
   371 => (x"97",x"cc",x"e5",x"c2"),
   372 => (x"d5",x"c1",x"49",x"bf"),
   373 => (x"cd",x"c0",x"05",x"a9"),
   374 => (x"cd",x"e5",x"c2",x"87"),
   375 => (x"c2",x"49",x"bf",x"97"),
   376 => (x"c0",x"02",x"a9",x"ea"),
   377 => (x"48",x"c0",x"87",x"c5"),
   378 => (x"c2",x"87",x"c7",x"c6"),
   379 => (x"bf",x"97",x"ce",x"dd"),
   380 => (x"e9",x"c3",x"48",x"7e"),
   381 => (x"ce",x"c0",x"02",x"a8"),
   382 => (x"c3",x"48",x"6e",x"87"),
   383 => (x"c0",x"02",x"a8",x"eb"),
   384 => (x"48",x"c0",x"87",x"c5"),
   385 => (x"c2",x"87",x"eb",x"c5"),
   386 => (x"bf",x"97",x"d9",x"dd"),
   387 => (x"c0",x"05",x"99",x"49"),
   388 => (x"dd",x"c2",x"87",x"cc"),
   389 => (x"49",x"bf",x"97",x"da"),
   390 => (x"c0",x"02",x"a9",x"c2"),
   391 => (x"48",x"c0",x"87",x"c5"),
   392 => (x"c2",x"87",x"cf",x"c5"),
   393 => (x"bf",x"97",x"db",x"dd"),
   394 => (x"d2",x"e5",x"c2",x"48"),
   395 => (x"48",x"4c",x"70",x"58"),
   396 => (x"e5",x"c2",x"88",x"c1"),
   397 => (x"dd",x"c2",x"58",x"d6"),
   398 => (x"49",x"bf",x"97",x"dc"),
   399 => (x"dd",x"c2",x"81",x"75"),
   400 => (x"4a",x"bf",x"97",x"dd"),
   401 => (x"a1",x"72",x"32",x"c8"),
   402 => (x"e3",x"e9",x"c2",x"7e"),
   403 => (x"c2",x"78",x"6e",x"48"),
   404 => (x"bf",x"97",x"de",x"dd"),
   405 => (x"58",x"a6",x"c8",x"48"),
   406 => (x"bf",x"d6",x"e5",x"c2"),
   407 => (x"87",x"d4",x"c2",x"02"),
   408 => (x"bf",x"c7",x"f2",x"c0"),
   409 => (x"e0",x"de",x"c2",x"49"),
   410 => (x"4b",x"c8",x"71",x"4a"),
   411 => (x"70",x"87",x"fb",x"e7"),
   412 => (x"c5",x"c0",x"02",x"98"),
   413 => (x"c3",x"48",x"c0",x"87"),
   414 => (x"e5",x"c2",x"87",x"f8"),
   415 => (x"c2",x"4c",x"bf",x"ce"),
   416 => (x"c2",x"5c",x"f7",x"e9"),
   417 => (x"bf",x"97",x"f3",x"dd"),
   418 => (x"c2",x"31",x"c8",x"49"),
   419 => (x"bf",x"97",x"f2",x"dd"),
   420 => (x"c2",x"49",x"a1",x"4a"),
   421 => (x"bf",x"97",x"f4",x"dd"),
   422 => (x"72",x"32",x"d0",x"4a"),
   423 => (x"dd",x"c2",x"49",x"a1"),
   424 => (x"4a",x"bf",x"97",x"f5"),
   425 => (x"a1",x"72",x"32",x"d8"),
   426 => (x"91",x"66",x"c4",x"49"),
   427 => (x"bf",x"e3",x"e9",x"c2"),
   428 => (x"eb",x"e9",x"c2",x"81"),
   429 => (x"fb",x"dd",x"c2",x"59"),
   430 => (x"c8",x"4a",x"bf",x"97"),
   431 => (x"fa",x"dd",x"c2",x"32"),
   432 => (x"a2",x"4b",x"bf",x"97"),
   433 => (x"fc",x"dd",x"c2",x"4a"),
   434 => (x"d0",x"4b",x"bf",x"97"),
   435 => (x"4a",x"a2",x"73",x"33"),
   436 => (x"97",x"fd",x"dd",x"c2"),
   437 => (x"9b",x"cf",x"4b",x"bf"),
   438 => (x"a2",x"73",x"33",x"d8"),
   439 => (x"ef",x"e9",x"c2",x"4a"),
   440 => (x"eb",x"e9",x"c2",x"5a"),
   441 => (x"8a",x"c2",x"4a",x"bf"),
   442 => (x"e9",x"c2",x"92",x"74"),
   443 => (x"a1",x"72",x"48",x"ef"),
   444 => (x"87",x"ca",x"c1",x"78"),
   445 => (x"97",x"e0",x"dd",x"c2"),
   446 => (x"31",x"c8",x"49",x"bf"),
   447 => (x"97",x"df",x"dd",x"c2"),
   448 => (x"49",x"a1",x"4a",x"bf"),
   449 => (x"59",x"de",x"e5",x"c2"),
   450 => (x"bf",x"da",x"e5",x"c2"),
   451 => (x"c7",x"31",x"c5",x"49"),
   452 => (x"29",x"c9",x"81",x"ff"),
   453 => (x"59",x"f7",x"e9",x"c2"),
   454 => (x"97",x"e5",x"dd",x"c2"),
   455 => (x"32",x"c8",x"4a",x"bf"),
   456 => (x"97",x"e4",x"dd",x"c2"),
   457 => (x"4a",x"a2",x"4b",x"bf"),
   458 => (x"6e",x"92",x"66",x"c4"),
   459 => (x"f3",x"e9",x"c2",x"82"),
   460 => (x"eb",x"e9",x"c2",x"5a"),
   461 => (x"c2",x"78",x"c0",x"48"),
   462 => (x"72",x"48",x"e7",x"e9"),
   463 => (x"e9",x"c2",x"78",x"a1"),
   464 => (x"e9",x"c2",x"48",x"f7"),
   465 => (x"c2",x"78",x"bf",x"eb"),
   466 => (x"c2",x"48",x"fb",x"e9"),
   467 => (x"78",x"bf",x"ef",x"e9"),
   468 => (x"bf",x"d6",x"e5",x"c2"),
   469 => (x"87",x"c9",x"c0",x"02"),
   470 => (x"30",x"c4",x"48",x"74"),
   471 => (x"c9",x"c0",x"7e",x"70"),
   472 => (x"f3",x"e9",x"c2",x"87"),
   473 => (x"30",x"c4",x"48",x"bf"),
   474 => (x"e5",x"c2",x"7e",x"70"),
   475 => (x"78",x"6e",x"48",x"da"),
   476 => (x"8e",x"f8",x"48",x"c1"),
   477 => (x"4c",x"26",x"4d",x"26"),
   478 => (x"4f",x"26",x"4b",x"26"),
   479 => (x"5c",x"5b",x"5e",x"0e"),
   480 => (x"4a",x"71",x"0e",x"5d"),
   481 => (x"bf",x"d6",x"e5",x"c2"),
   482 => (x"72",x"87",x"cb",x"02"),
   483 => (x"72",x"2b",x"c7",x"4b"),
   484 => (x"9c",x"ff",x"c1",x"4c"),
   485 => (x"4b",x"72",x"87",x"c9"),
   486 => (x"4c",x"72",x"2b",x"c8"),
   487 => (x"c2",x"9c",x"ff",x"c3"),
   488 => (x"83",x"bf",x"e3",x"e9"),
   489 => (x"bf",x"c3",x"f2",x"c0"),
   490 => (x"87",x"d9",x"02",x"ab"),
   491 => (x"5b",x"c7",x"f2",x"c0"),
   492 => (x"1e",x"ce",x"dd",x"c2"),
   493 => (x"fd",x"f0",x"49",x"73"),
   494 => (x"70",x"86",x"c4",x"87"),
   495 => (x"87",x"c5",x"05",x"98"),
   496 => (x"e6",x"c0",x"48",x"c0"),
   497 => (x"d6",x"e5",x"c2",x"87"),
   498 => (x"87",x"d2",x"02",x"bf"),
   499 => (x"91",x"c4",x"49",x"74"),
   500 => (x"81",x"ce",x"dd",x"c2"),
   501 => (x"ff",x"cf",x"4d",x"69"),
   502 => (x"9d",x"ff",x"ff",x"ff"),
   503 => (x"49",x"74",x"87",x"cb"),
   504 => (x"dd",x"c2",x"91",x"c2"),
   505 => (x"69",x"9f",x"81",x"ce"),
   506 => (x"fe",x"48",x"75",x"4d"),
   507 => (x"5e",x"0e",x"87",x"c6"),
   508 => (x"0e",x"5d",x"5c",x"5b"),
   509 => (x"c0",x"4d",x"71",x"1e"),
   510 => (x"ca",x"49",x"c1",x"1e"),
   511 => (x"86",x"c4",x"87",x"ee"),
   512 => (x"02",x"9c",x"4c",x"70"),
   513 => (x"c2",x"87",x"c0",x"c1"),
   514 => (x"75",x"4a",x"de",x"e5"),
   515 => (x"87",x"ff",x"e0",x"49"),
   516 => (x"c0",x"02",x"98",x"70"),
   517 => (x"4a",x"74",x"87",x"f1"),
   518 => (x"4b",x"cb",x"49",x"75"),
   519 => (x"70",x"87",x"e5",x"e1"),
   520 => (x"e2",x"c0",x"02",x"98"),
   521 => (x"74",x"1e",x"c0",x"87"),
   522 => (x"87",x"c7",x"02",x"9c"),
   523 => (x"c0",x"48",x"a6",x"c4"),
   524 => (x"c4",x"87",x"c5",x"78"),
   525 => (x"78",x"c1",x"48",x"a6"),
   526 => (x"c9",x"49",x"66",x"c4"),
   527 => (x"86",x"c4",x"87",x"ee"),
   528 => (x"05",x"9c",x"4c",x"70"),
   529 => (x"74",x"87",x"c0",x"ff"),
   530 => (x"e7",x"fc",x"26",x"48"),
   531 => (x"5b",x"5e",x"0e",x"87"),
   532 => (x"1e",x"0e",x"5d",x"5c"),
   533 => (x"05",x"9b",x"4b",x"71"),
   534 => (x"48",x"c0",x"87",x"c5"),
   535 => (x"c8",x"87",x"e5",x"c1"),
   536 => (x"7d",x"c0",x"4d",x"a3"),
   537 => (x"c7",x"02",x"66",x"d4"),
   538 => (x"97",x"66",x"d4",x"87"),
   539 => (x"87",x"c5",x"05",x"bf"),
   540 => (x"cf",x"c1",x"48",x"c0"),
   541 => (x"49",x"66",x"d4",x"87"),
   542 => (x"70",x"87",x"f3",x"fd"),
   543 => (x"c1",x"02",x"9c",x"4c"),
   544 => (x"a4",x"dc",x"87",x"c0"),
   545 => (x"da",x"7d",x"69",x"49"),
   546 => (x"a3",x"c4",x"49",x"a4"),
   547 => (x"7a",x"69",x"9f",x"4a"),
   548 => (x"bf",x"d6",x"e5",x"c2"),
   549 => (x"d4",x"87",x"d2",x"02"),
   550 => (x"69",x"9f",x"49",x"a4"),
   551 => (x"ff",x"ff",x"c0",x"49"),
   552 => (x"d0",x"48",x"71",x"99"),
   553 => (x"c2",x"7e",x"70",x"30"),
   554 => (x"6e",x"7e",x"c0",x"87"),
   555 => (x"80",x"6a",x"48",x"49"),
   556 => (x"7b",x"c0",x"7a",x"70"),
   557 => (x"6a",x"49",x"a3",x"cc"),
   558 => (x"49",x"a3",x"d0",x"79"),
   559 => (x"48",x"74",x"79",x"c0"),
   560 => (x"48",x"c0",x"87",x"c2"),
   561 => (x"87",x"ec",x"fa",x"26"),
   562 => (x"5c",x"5b",x"5e",x"0e"),
   563 => (x"4c",x"71",x"0e",x"5d"),
   564 => (x"48",x"c3",x"f2",x"c0"),
   565 => (x"9c",x"74",x"78",x"ff"),
   566 => (x"87",x"ca",x"c1",x"02"),
   567 => (x"69",x"49",x"a4",x"c8"),
   568 => (x"87",x"c2",x"c1",x"02"),
   569 => (x"6c",x"4a",x"66",x"d0"),
   570 => (x"a6",x"d4",x"82",x"49"),
   571 => (x"4d",x"66",x"d0",x"5a"),
   572 => (x"d2",x"e5",x"c2",x"b9"),
   573 => (x"ba",x"ff",x"4a",x"bf"),
   574 => (x"99",x"71",x"99",x"72"),
   575 => (x"87",x"e4",x"c0",x"02"),
   576 => (x"6b",x"4b",x"a4",x"c4"),
   577 => (x"87",x"f4",x"f9",x"49"),
   578 => (x"e5",x"c2",x"7b",x"70"),
   579 => (x"6c",x"49",x"bf",x"ce"),
   580 => (x"75",x"7c",x"71",x"81"),
   581 => (x"d2",x"e5",x"c2",x"b9"),
   582 => (x"ba",x"ff",x"4a",x"bf"),
   583 => (x"99",x"71",x"99",x"72"),
   584 => (x"87",x"dc",x"ff",x"05"),
   585 => (x"cb",x"f9",x"7c",x"75"),
   586 => (x"1e",x"73",x"1e",x"87"),
   587 => (x"02",x"9b",x"4b",x"71"),
   588 => (x"a3",x"c8",x"87",x"c7"),
   589 => (x"c5",x"05",x"69",x"49"),
   590 => (x"c0",x"48",x"c0",x"87"),
   591 => (x"e9",x"c2",x"87",x"eb"),
   592 => (x"c4",x"4a",x"bf",x"e7"),
   593 => (x"49",x"69",x"49",x"a3"),
   594 => (x"e5",x"c2",x"89",x"c2"),
   595 => (x"71",x"91",x"bf",x"ce"),
   596 => (x"e5",x"c2",x"4a",x"a2"),
   597 => (x"6b",x"49",x"bf",x"d2"),
   598 => (x"4a",x"a2",x"71",x"99"),
   599 => (x"72",x"1e",x"66",x"c8"),
   600 => (x"87",x"d2",x"ea",x"49"),
   601 => (x"49",x"70",x"86",x"c4"),
   602 => (x"87",x"cc",x"f8",x"48"),
   603 => (x"71",x"1e",x"73",x"1e"),
   604 => (x"c7",x"02",x"9b",x"4b"),
   605 => (x"49",x"a3",x"c8",x"87"),
   606 => (x"87",x"c5",x"05",x"69"),
   607 => (x"eb",x"c0",x"48",x"c0"),
   608 => (x"e7",x"e9",x"c2",x"87"),
   609 => (x"a3",x"c4",x"4a",x"bf"),
   610 => (x"c2",x"49",x"69",x"49"),
   611 => (x"ce",x"e5",x"c2",x"89"),
   612 => (x"a2",x"71",x"91",x"bf"),
   613 => (x"d2",x"e5",x"c2",x"4a"),
   614 => (x"99",x"6b",x"49",x"bf"),
   615 => (x"c8",x"4a",x"a2",x"71"),
   616 => (x"49",x"72",x"1e",x"66"),
   617 => (x"c4",x"87",x"c5",x"e6"),
   618 => (x"48",x"49",x"70",x"86"),
   619 => (x"0e",x"87",x"c9",x"f7"),
   620 => (x"5d",x"5c",x"5b",x"5e"),
   621 => (x"4b",x"71",x"1e",x"0e"),
   622 => (x"c9",x"4c",x"66",x"d4"),
   623 => (x"02",x"9b",x"73",x"2c"),
   624 => (x"c8",x"87",x"cf",x"c1"),
   625 => (x"02",x"69",x"49",x"a3"),
   626 => (x"d0",x"87",x"c7",x"c1"),
   627 => (x"66",x"d4",x"4d",x"a3"),
   628 => (x"d2",x"e5",x"c2",x"7d"),
   629 => (x"b9",x"ff",x"49",x"bf"),
   630 => (x"7e",x"99",x"4a",x"6b"),
   631 => (x"cd",x"03",x"ac",x"71"),
   632 => (x"7d",x"7b",x"c0",x"87"),
   633 => (x"c4",x"4a",x"a3",x"cc"),
   634 => (x"79",x"6a",x"49",x"a3"),
   635 => (x"8c",x"72",x"87",x"c2"),
   636 => (x"dd",x"02",x"9c",x"74"),
   637 => (x"73",x"1e",x"49",x"87"),
   638 => (x"87",x"cc",x"fb",x"49"),
   639 => (x"66",x"d4",x"86",x"c4"),
   640 => (x"99",x"ff",x"c7",x"49"),
   641 => (x"c2",x"87",x"cb",x"02"),
   642 => (x"73",x"1e",x"ce",x"dd"),
   643 => (x"87",x"d9",x"fc",x"49"),
   644 => (x"f5",x"26",x"86",x"c4"),
   645 => (x"73",x"1e",x"87",x"de"),
   646 => (x"9b",x"4b",x"71",x"1e"),
   647 => (x"87",x"e4",x"c0",x"02"),
   648 => (x"5b",x"fb",x"e9",x"c2"),
   649 => (x"8a",x"c2",x"4a",x"73"),
   650 => (x"bf",x"ce",x"e5",x"c2"),
   651 => (x"e9",x"c2",x"92",x"49"),
   652 => (x"72",x"48",x"bf",x"e7"),
   653 => (x"ff",x"e9",x"c2",x"80"),
   654 => (x"c4",x"48",x"71",x"58"),
   655 => (x"de",x"e5",x"c2",x"30"),
   656 => (x"87",x"ed",x"c0",x"58"),
   657 => (x"48",x"f7",x"e9",x"c2"),
   658 => (x"bf",x"eb",x"e9",x"c2"),
   659 => (x"fb",x"e9",x"c2",x"78"),
   660 => (x"ef",x"e9",x"c2",x"48"),
   661 => (x"e5",x"c2",x"78",x"bf"),
   662 => (x"c9",x"02",x"bf",x"d6"),
   663 => (x"ce",x"e5",x"c2",x"87"),
   664 => (x"31",x"c4",x"49",x"bf"),
   665 => (x"e9",x"c2",x"87",x"c7"),
   666 => (x"c4",x"49",x"bf",x"f3"),
   667 => (x"de",x"e5",x"c2",x"31"),
   668 => (x"87",x"c4",x"f4",x"59"),
   669 => (x"5c",x"5b",x"5e",x"0e"),
   670 => (x"c0",x"4a",x"71",x"0e"),
   671 => (x"02",x"9a",x"72",x"4b"),
   672 => (x"da",x"87",x"e1",x"c0"),
   673 => (x"69",x"9f",x"49",x"a2"),
   674 => (x"d6",x"e5",x"c2",x"4b"),
   675 => (x"87",x"cf",x"02",x"bf"),
   676 => (x"9f",x"49",x"a2",x"d4"),
   677 => (x"c0",x"4c",x"49",x"69"),
   678 => (x"d0",x"9c",x"ff",x"ff"),
   679 => (x"c0",x"87",x"c2",x"34"),
   680 => (x"b3",x"49",x"74",x"4c"),
   681 => (x"ed",x"fd",x"49",x"73"),
   682 => (x"87",x"ca",x"f3",x"87"),
   683 => (x"5c",x"5b",x"5e",x"0e"),
   684 => (x"86",x"f4",x"0e",x"5d"),
   685 => (x"7e",x"c0",x"4a",x"71"),
   686 => (x"d8",x"02",x"9a",x"72"),
   687 => (x"ca",x"dd",x"c2",x"87"),
   688 => (x"c2",x"78",x"c0",x"48"),
   689 => (x"c2",x"48",x"c2",x"dd"),
   690 => (x"78",x"bf",x"fb",x"e9"),
   691 => (x"48",x"c6",x"dd",x"c2"),
   692 => (x"bf",x"f7",x"e9",x"c2"),
   693 => (x"eb",x"e5",x"c2",x"78"),
   694 => (x"c2",x"50",x"c0",x"48"),
   695 => (x"49",x"bf",x"da",x"e5"),
   696 => (x"bf",x"ca",x"dd",x"c2"),
   697 => (x"03",x"aa",x"71",x"4a"),
   698 => (x"72",x"87",x"ff",x"c3"),
   699 => (x"05",x"99",x"cf",x"49"),
   700 => (x"c2",x"87",x"e0",x"c0"),
   701 => (x"c2",x"1e",x"ce",x"dd"),
   702 => (x"49",x"bf",x"c2",x"dd"),
   703 => (x"48",x"c2",x"dd",x"c2"),
   704 => (x"71",x"78",x"a1",x"c1"),
   705 => (x"c4",x"87",x"ef",x"e3"),
   706 => (x"ff",x"f1",x"c0",x"86"),
   707 => (x"ce",x"dd",x"c2",x"48"),
   708 => (x"c0",x"87",x"cc",x"78"),
   709 => (x"48",x"bf",x"ff",x"f1"),
   710 => (x"c0",x"80",x"e0",x"c0"),
   711 => (x"c2",x"58",x"c3",x"f2"),
   712 => (x"48",x"bf",x"ca",x"dd"),
   713 => (x"dd",x"c2",x"80",x"c1"),
   714 => (x"7f",x"27",x"58",x"ce"),
   715 => (x"bf",x"00",x"00",x"0c"),
   716 => (x"9d",x"4d",x"bf",x"97"),
   717 => (x"87",x"e2",x"c2",x"02"),
   718 => (x"02",x"ad",x"e5",x"c3"),
   719 => (x"c0",x"87",x"db",x"c2"),
   720 => (x"4b",x"bf",x"ff",x"f1"),
   721 => (x"11",x"49",x"a3",x"cb"),
   722 => (x"05",x"ac",x"cf",x"4c"),
   723 => (x"75",x"87",x"d2",x"c1"),
   724 => (x"c1",x"99",x"df",x"49"),
   725 => (x"c2",x"91",x"cd",x"89"),
   726 => (x"c1",x"81",x"de",x"e5"),
   727 => (x"51",x"12",x"4a",x"a3"),
   728 => (x"12",x"4a",x"a3",x"c3"),
   729 => (x"4a",x"a3",x"c5",x"51"),
   730 => (x"a3",x"c7",x"51",x"12"),
   731 => (x"c9",x"51",x"12",x"4a"),
   732 => (x"51",x"12",x"4a",x"a3"),
   733 => (x"12",x"4a",x"a3",x"ce"),
   734 => (x"4a",x"a3",x"d0",x"51"),
   735 => (x"a3",x"d2",x"51",x"12"),
   736 => (x"d4",x"51",x"12",x"4a"),
   737 => (x"51",x"12",x"4a",x"a3"),
   738 => (x"12",x"4a",x"a3",x"d6"),
   739 => (x"4a",x"a3",x"d8",x"51"),
   740 => (x"a3",x"dc",x"51",x"12"),
   741 => (x"de",x"51",x"12",x"4a"),
   742 => (x"51",x"12",x"4a",x"a3"),
   743 => (x"f9",x"c0",x"7e",x"c1"),
   744 => (x"c8",x"49",x"74",x"87"),
   745 => (x"ea",x"c0",x"05",x"99"),
   746 => (x"d0",x"49",x"74",x"87"),
   747 => (x"87",x"d0",x"05",x"99"),
   748 => (x"c0",x"02",x"66",x"dc"),
   749 => (x"49",x"73",x"87",x"ca"),
   750 => (x"70",x"0f",x"66",x"dc"),
   751 => (x"87",x"d3",x"02",x"98"),
   752 => (x"c6",x"c0",x"05",x"6e"),
   753 => (x"de",x"e5",x"c2",x"87"),
   754 => (x"c0",x"50",x"c0",x"48"),
   755 => (x"48",x"bf",x"ff",x"f1"),
   756 => (x"c2",x"87",x"e7",x"c2"),
   757 => (x"c0",x"48",x"eb",x"e5"),
   758 => (x"e5",x"c2",x"7e",x"50"),
   759 => (x"c2",x"49",x"bf",x"da"),
   760 => (x"4a",x"bf",x"ca",x"dd"),
   761 => (x"fc",x"04",x"aa",x"71"),
   762 => (x"e9",x"c2",x"87",x"c1"),
   763 => (x"c0",x"05",x"bf",x"fb"),
   764 => (x"e5",x"c2",x"87",x"c8"),
   765 => (x"c1",x"02",x"bf",x"d6"),
   766 => (x"f2",x"c0",x"87",x"fe"),
   767 => (x"78",x"ff",x"48",x"c3"),
   768 => (x"bf",x"c6",x"dd",x"c2"),
   769 => (x"87",x"f4",x"ed",x"49"),
   770 => (x"dd",x"c2",x"49",x"70"),
   771 => (x"a6",x"c4",x"59",x"ca"),
   772 => (x"c6",x"dd",x"c2",x"48"),
   773 => (x"e5",x"c2",x"78",x"bf"),
   774 => (x"c0",x"02",x"bf",x"d6"),
   775 => (x"66",x"c4",x"87",x"d8"),
   776 => (x"ff",x"ff",x"cf",x"49"),
   777 => (x"a9",x"99",x"f8",x"ff"),
   778 => (x"87",x"c5",x"c0",x"02"),
   779 => (x"e1",x"c0",x"4d",x"c0"),
   780 => (x"c0",x"4d",x"c1",x"87"),
   781 => (x"66",x"c4",x"87",x"dc"),
   782 => (x"f8",x"ff",x"cf",x"49"),
   783 => (x"c0",x"02",x"a9",x"99"),
   784 => (x"a6",x"c8",x"87",x"c8"),
   785 => (x"c0",x"78",x"c0",x"48"),
   786 => (x"a6",x"c8",x"87",x"c5"),
   787 => (x"c8",x"78",x"c1",x"48"),
   788 => (x"9d",x"75",x"4d",x"66"),
   789 => (x"87",x"e0",x"c0",x"05"),
   790 => (x"c2",x"49",x"66",x"c4"),
   791 => (x"ce",x"e5",x"c2",x"89"),
   792 => (x"c2",x"91",x"4a",x"bf"),
   793 => (x"4a",x"bf",x"e7",x"e9"),
   794 => (x"48",x"c2",x"dd",x"c2"),
   795 => (x"c2",x"78",x"a1",x"72"),
   796 => (x"c0",x"48",x"ca",x"dd"),
   797 => (x"87",x"e3",x"f9",x"78"),
   798 => (x"8e",x"f4",x"48",x"c0"),
   799 => (x"00",x"87",x"f5",x"eb"),
   800 => (x"ff",x"00",x"00",x"00"),
   801 => (x"8f",x"ff",x"ff",x"ff"),
   802 => (x"98",x"00",x"00",x"0c"),
   803 => (x"46",x"00",x"00",x"0c"),
   804 => (x"32",x"33",x"54",x"41"),
   805 => (x"00",x"20",x"20",x"20"),
   806 => (x"31",x"54",x"41",x"46"),
   807 => (x"20",x"20",x"20",x"36"),
   808 => (x"d4",x"ff",x"1e",x"00"),
   809 => (x"78",x"ff",x"c3",x"48"),
   810 => (x"4f",x"26",x"48",x"68"),
   811 => (x"48",x"d4",x"ff",x"1e"),
   812 => (x"ff",x"78",x"ff",x"c3"),
   813 => (x"e1",x"c8",x"48",x"d0"),
   814 => (x"48",x"d4",x"ff",x"78"),
   815 => (x"e9",x"c2",x"78",x"d4"),
   816 => (x"d4",x"ff",x"48",x"ff"),
   817 => (x"4f",x"26",x"50",x"bf"),
   818 => (x"48",x"d0",x"ff",x"1e"),
   819 => (x"26",x"78",x"e0",x"c0"),
   820 => (x"cc",x"ff",x"1e",x"4f"),
   821 => (x"99",x"49",x"70",x"87"),
   822 => (x"c0",x"87",x"c6",x"02"),
   823 => (x"f1",x"05",x"a9",x"fb"),
   824 => (x"26",x"48",x"71",x"87"),
   825 => (x"5b",x"5e",x"0e",x"4f"),
   826 => (x"4b",x"71",x"0e",x"5c"),
   827 => (x"f0",x"fe",x"4c",x"c0"),
   828 => (x"99",x"49",x"70",x"87"),
   829 => (x"87",x"f9",x"c0",x"02"),
   830 => (x"02",x"a9",x"ec",x"c0"),
   831 => (x"c0",x"87",x"f2",x"c0"),
   832 => (x"c0",x"02",x"a9",x"fb"),
   833 => (x"66",x"cc",x"87",x"eb"),
   834 => (x"c7",x"03",x"ac",x"b7"),
   835 => (x"02",x"66",x"d0",x"87"),
   836 => (x"53",x"71",x"87",x"c2"),
   837 => (x"c2",x"02",x"99",x"71"),
   838 => (x"fe",x"84",x"c1",x"87"),
   839 => (x"49",x"70",x"87",x"c3"),
   840 => (x"87",x"cd",x"02",x"99"),
   841 => (x"02",x"a9",x"ec",x"c0"),
   842 => (x"fb",x"c0",x"87",x"c7"),
   843 => (x"d5",x"ff",x"05",x"a9"),
   844 => (x"02",x"66",x"d0",x"87"),
   845 => (x"97",x"c0",x"87",x"c3"),
   846 => (x"a9",x"ec",x"c0",x"7b"),
   847 => (x"74",x"87",x"c4",x"05"),
   848 => (x"74",x"87",x"c5",x"4a"),
   849 => (x"8a",x"0a",x"c0",x"4a"),
   850 => (x"87",x"c2",x"48",x"72"),
   851 => (x"4c",x"26",x"4d",x"26"),
   852 => (x"4f",x"26",x"4b",x"26"),
   853 => (x"87",x"c9",x"fd",x"1e"),
   854 => (x"f0",x"c0",x"49",x"70"),
   855 => (x"ca",x"04",x"a9",x"b7"),
   856 => (x"b7",x"f9",x"c0",x"87"),
   857 => (x"87",x"c3",x"01",x"a9"),
   858 => (x"c1",x"89",x"f0",x"c0"),
   859 => (x"04",x"a9",x"b7",x"c1"),
   860 => (x"da",x"c1",x"87",x"ca"),
   861 => (x"c3",x"01",x"a9",x"b7"),
   862 => (x"89",x"f7",x"c0",x"87"),
   863 => (x"4f",x"26",x"48",x"71"),
   864 => (x"5c",x"5b",x"5e",x"0e"),
   865 => (x"ff",x"4a",x"71",x"0e"),
   866 => (x"49",x"72",x"4c",x"d4"),
   867 => (x"70",x"87",x"ea",x"c0"),
   868 => (x"c2",x"02",x"9b",x"4b"),
   869 => (x"ff",x"8b",x"c1",x"87"),
   870 => (x"c5",x"c8",x"48",x"d0"),
   871 => (x"7c",x"d5",x"c1",x"78"),
   872 => (x"31",x"c6",x"49",x"73"),
   873 => (x"97",x"d2",x"db",x"c2"),
   874 => (x"71",x"48",x"4a",x"bf"),
   875 => (x"ff",x"7c",x"70",x"b0"),
   876 => (x"78",x"c4",x"48",x"d0"),
   877 => (x"d5",x"fe",x"48",x"73"),
   878 => (x"5b",x"5e",x"0e",x"87"),
   879 => (x"f8",x"0e",x"5d",x"5c"),
   880 => (x"c0",x"4c",x"71",x"86"),
   881 => (x"87",x"e4",x"fb",x"7e"),
   882 => (x"f9",x"c0",x"4b",x"c0"),
   883 => (x"49",x"bf",x"97",x"e6"),
   884 => (x"cf",x"04",x"a9",x"c0"),
   885 => (x"87",x"f9",x"fb",x"87"),
   886 => (x"f9",x"c0",x"83",x"c1"),
   887 => (x"49",x"bf",x"97",x"e6"),
   888 => (x"87",x"f1",x"06",x"ab"),
   889 => (x"97",x"e6",x"f9",x"c0"),
   890 => (x"87",x"cf",x"02",x"bf"),
   891 => (x"70",x"87",x"f2",x"fa"),
   892 => (x"c6",x"02",x"99",x"49"),
   893 => (x"a9",x"ec",x"c0",x"87"),
   894 => (x"c0",x"87",x"f1",x"05"),
   895 => (x"87",x"e1",x"fa",x"4b"),
   896 => (x"dc",x"fa",x"4d",x"70"),
   897 => (x"58",x"a6",x"c8",x"87"),
   898 => (x"70",x"87",x"d6",x"fa"),
   899 => (x"c8",x"83",x"c1",x"4a"),
   900 => (x"69",x"97",x"49",x"a4"),
   901 => (x"c7",x"02",x"ad",x"49"),
   902 => (x"ad",x"ff",x"c0",x"87"),
   903 => (x"87",x"e7",x"c0",x"05"),
   904 => (x"97",x"49",x"a4",x"c9"),
   905 => (x"66",x"c4",x"49",x"69"),
   906 => (x"87",x"c7",x"02",x"a9"),
   907 => (x"a8",x"ff",x"c0",x"48"),
   908 => (x"ca",x"87",x"d4",x"05"),
   909 => (x"69",x"97",x"49",x"a4"),
   910 => (x"c6",x"02",x"aa",x"49"),
   911 => (x"aa",x"ff",x"c0",x"87"),
   912 => (x"c1",x"87",x"c4",x"05"),
   913 => (x"c0",x"87",x"d0",x"7e"),
   914 => (x"c6",x"02",x"ad",x"ec"),
   915 => (x"ad",x"fb",x"c0",x"87"),
   916 => (x"c0",x"87",x"c4",x"05"),
   917 => (x"6e",x"7e",x"c1",x"4b"),
   918 => (x"87",x"e1",x"fe",x"02"),
   919 => (x"73",x"87",x"e9",x"f9"),
   920 => (x"fb",x"8e",x"f8",x"48"),
   921 => (x"0e",x"00",x"87",x"e6"),
   922 => (x"5d",x"5c",x"5b",x"5e"),
   923 => (x"4b",x"71",x"1e",x"0e"),
   924 => (x"ab",x"4d",x"4c",x"c0"),
   925 => (x"87",x"e8",x"c0",x"04"),
   926 => (x"1e",x"f9",x"f6",x"c0"),
   927 => (x"c4",x"02",x"9d",x"75"),
   928 => (x"c2",x"4a",x"c0",x"87"),
   929 => (x"72",x"4a",x"c1",x"87"),
   930 => (x"87",x"e0",x"f0",x"49"),
   931 => (x"7e",x"70",x"86",x"c4"),
   932 => (x"05",x"6e",x"84",x"c1"),
   933 => (x"4c",x"73",x"87",x"c2"),
   934 => (x"ac",x"73",x"85",x"c1"),
   935 => (x"87",x"d8",x"ff",x"06"),
   936 => (x"26",x"26",x"48",x"6e"),
   937 => (x"26",x"4c",x"26",x"4d"),
   938 => (x"0e",x"4f",x"26",x"4b"),
   939 => (x"5d",x"5c",x"5b",x"5e"),
   940 => (x"4c",x"71",x"1e",x"0e"),
   941 => (x"c2",x"91",x"de",x"49"),
   942 => (x"71",x"4d",x"d9",x"ea"),
   943 => (x"02",x"6d",x"97",x"85"),
   944 => (x"c2",x"87",x"dd",x"c1"),
   945 => (x"4a",x"bf",x"c4",x"ea"),
   946 => (x"49",x"72",x"82",x"74"),
   947 => (x"70",x"87",x"d8",x"fe"),
   948 => (x"c0",x"02",x"6e",x"7e"),
   949 => (x"ea",x"c2",x"87",x"f3"),
   950 => (x"4a",x"6e",x"4b",x"cc"),
   951 => (x"c7",x"ff",x"49",x"cb"),
   952 => (x"4b",x"74",x"87",x"c6"),
   953 => (x"dd",x"c1",x"93",x"cb"),
   954 => (x"83",x"c4",x"83",x"fa"),
   955 => (x"7b",x"e4",x"fc",x"c0"),
   956 => (x"c3",x"c1",x"49",x"74"),
   957 => (x"7b",x"75",x"87",x"f3"),
   958 => (x"97",x"d8",x"ea",x"c2"),
   959 => (x"c2",x"1e",x"49",x"bf"),
   960 => (x"c1",x"49",x"cc",x"ea"),
   961 => (x"c4",x"87",x"cd",x"de"),
   962 => (x"c1",x"49",x"74",x"86"),
   963 => (x"c0",x"87",x"da",x"c3"),
   964 => (x"f9",x"c4",x"c1",x"49"),
   965 => (x"c0",x"ea",x"c2",x"87"),
   966 => (x"c1",x"78",x"c0",x"48"),
   967 => (x"87",x"cb",x"dd",x"49"),
   968 => (x"87",x"ff",x"fd",x"26"),
   969 => (x"64",x"61",x"6f",x"4c"),
   970 => (x"2e",x"67",x"6e",x"69"),
   971 => (x"0e",x"00",x"2e",x"2e"),
   972 => (x"0e",x"5c",x"5b",x"5e"),
   973 => (x"c2",x"4a",x"4b",x"71"),
   974 => (x"82",x"bf",x"c4",x"ea"),
   975 => (x"e6",x"fc",x"49",x"72"),
   976 => (x"9c",x"4c",x"70",x"87"),
   977 => (x"49",x"87",x"c4",x"02"),
   978 => (x"c2",x"87",x"e9",x"ec"),
   979 => (x"c0",x"48",x"c4",x"ea"),
   980 => (x"dc",x"49",x"c1",x"78"),
   981 => (x"cc",x"fd",x"87",x"d5"),
   982 => (x"5b",x"5e",x"0e",x"87"),
   983 => (x"f4",x"0e",x"5d",x"5c"),
   984 => (x"ce",x"dd",x"c2",x"86"),
   985 => (x"c4",x"4c",x"c0",x"4d"),
   986 => (x"78",x"c0",x"48",x"a6"),
   987 => (x"bf",x"c4",x"ea",x"c2"),
   988 => (x"06",x"a9",x"c0",x"49"),
   989 => (x"c2",x"87",x"c1",x"c1"),
   990 => (x"98",x"48",x"ce",x"dd"),
   991 => (x"87",x"f8",x"c0",x"02"),
   992 => (x"1e",x"f9",x"f6",x"c0"),
   993 => (x"c7",x"02",x"66",x"c8"),
   994 => (x"48",x"a6",x"c4",x"87"),
   995 => (x"87",x"c5",x"78",x"c0"),
   996 => (x"c1",x"48",x"a6",x"c4"),
   997 => (x"49",x"66",x"c4",x"78"),
   998 => (x"c4",x"87",x"d1",x"ec"),
   999 => (x"c1",x"4d",x"70",x"86"),
  1000 => (x"48",x"66",x"c4",x"84"),
  1001 => (x"a6",x"c8",x"80",x"c1"),
  1002 => (x"c4",x"ea",x"c2",x"58"),
  1003 => (x"03",x"ac",x"49",x"bf"),
  1004 => (x"9d",x"75",x"87",x"c6"),
  1005 => (x"87",x"c8",x"ff",x"05"),
  1006 => (x"9d",x"75",x"4c",x"c0"),
  1007 => (x"87",x"e0",x"c3",x"02"),
  1008 => (x"1e",x"f9",x"f6",x"c0"),
  1009 => (x"c7",x"02",x"66",x"c8"),
  1010 => (x"48",x"a6",x"cc",x"87"),
  1011 => (x"87",x"c5",x"78",x"c0"),
  1012 => (x"c1",x"48",x"a6",x"cc"),
  1013 => (x"49",x"66",x"cc",x"78"),
  1014 => (x"c4",x"87",x"d1",x"eb"),
  1015 => (x"6e",x"7e",x"70",x"86"),
  1016 => (x"87",x"e9",x"c2",x"02"),
  1017 => (x"81",x"cb",x"49",x"6e"),
  1018 => (x"d0",x"49",x"69",x"97"),
  1019 => (x"d6",x"c1",x"02",x"99"),
  1020 => (x"ef",x"fc",x"c0",x"87"),
  1021 => (x"cb",x"49",x"74",x"4a"),
  1022 => (x"fa",x"dd",x"c1",x"91"),
  1023 => (x"c8",x"79",x"72",x"81"),
  1024 => (x"51",x"ff",x"c3",x"81"),
  1025 => (x"91",x"de",x"49",x"74"),
  1026 => (x"4d",x"d9",x"ea",x"c2"),
  1027 => (x"c1",x"c2",x"85",x"71"),
  1028 => (x"a5",x"c1",x"7d",x"97"),
  1029 => (x"51",x"e0",x"c0",x"49"),
  1030 => (x"97",x"de",x"e5",x"c2"),
  1031 => (x"87",x"d2",x"02",x"bf"),
  1032 => (x"a5",x"c2",x"84",x"c1"),
  1033 => (x"de",x"e5",x"c2",x"4b"),
  1034 => (x"ff",x"49",x"db",x"4a"),
  1035 => (x"c1",x"87",x"f9",x"c1"),
  1036 => (x"a5",x"cd",x"87",x"db"),
  1037 => (x"c1",x"51",x"c0",x"49"),
  1038 => (x"4b",x"a5",x"c2",x"84"),
  1039 => (x"49",x"cb",x"4a",x"6e"),
  1040 => (x"87",x"e4",x"c1",x"ff"),
  1041 => (x"c0",x"87",x"c6",x"c1"),
  1042 => (x"74",x"4a",x"eb",x"fa"),
  1043 => (x"c1",x"91",x"cb",x"49"),
  1044 => (x"72",x"81",x"fa",x"dd"),
  1045 => (x"de",x"e5",x"c2",x"79"),
  1046 => (x"d8",x"02",x"bf",x"97"),
  1047 => (x"de",x"49",x"74",x"87"),
  1048 => (x"c2",x"84",x"c1",x"91"),
  1049 => (x"71",x"4b",x"d9",x"ea"),
  1050 => (x"de",x"e5",x"c2",x"83"),
  1051 => (x"ff",x"49",x"dd",x"4a"),
  1052 => (x"d8",x"87",x"f5",x"c0"),
  1053 => (x"de",x"4b",x"74",x"87"),
  1054 => (x"d9",x"ea",x"c2",x"93"),
  1055 => (x"49",x"a3",x"cb",x"83"),
  1056 => (x"84",x"c1",x"51",x"c0"),
  1057 => (x"cb",x"4a",x"6e",x"73"),
  1058 => (x"db",x"c0",x"ff",x"49"),
  1059 => (x"48",x"66",x"c4",x"87"),
  1060 => (x"a6",x"c8",x"80",x"c1"),
  1061 => (x"03",x"ac",x"c7",x"58"),
  1062 => (x"6e",x"87",x"c5",x"c0"),
  1063 => (x"87",x"e0",x"fc",x"05"),
  1064 => (x"8e",x"f4",x"48",x"74"),
  1065 => (x"1e",x"87",x"fc",x"f7"),
  1066 => (x"4b",x"71",x"1e",x"73"),
  1067 => (x"c1",x"91",x"cb",x"49"),
  1068 => (x"c8",x"81",x"fa",x"dd"),
  1069 => (x"db",x"c2",x"4a",x"a1"),
  1070 => (x"50",x"12",x"48",x"d2"),
  1071 => (x"c0",x"4a",x"a1",x"c9"),
  1072 => (x"12",x"48",x"e6",x"f9"),
  1073 => (x"c2",x"81",x"ca",x"50"),
  1074 => (x"11",x"48",x"d8",x"ea"),
  1075 => (x"d8",x"ea",x"c2",x"50"),
  1076 => (x"1e",x"49",x"bf",x"97"),
  1077 => (x"d6",x"c1",x"49",x"c0"),
  1078 => (x"ea",x"c2",x"87",x"fa"),
  1079 => (x"78",x"de",x"48",x"c0"),
  1080 => (x"c6",x"d6",x"49",x"c1"),
  1081 => (x"fe",x"f6",x"26",x"87"),
  1082 => (x"4a",x"71",x"1e",x"87"),
  1083 => (x"c1",x"91",x"cb",x"49"),
  1084 => (x"c8",x"81",x"fa",x"dd"),
  1085 => (x"c2",x"48",x"11",x"81"),
  1086 => (x"c2",x"58",x"c4",x"ea"),
  1087 => (x"c0",x"48",x"c4",x"ea"),
  1088 => (x"d5",x"49",x"c1",x"78"),
  1089 => (x"4f",x"26",x"87",x"e5"),
  1090 => (x"c0",x"49",x"c0",x"1e"),
  1091 => (x"26",x"87",x"ff",x"fc"),
  1092 => (x"99",x"71",x"1e",x"4f"),
  1093 => (x"c1",x"87",x"d2",x"02"),
  1094 => (x"c0",x"48",x"cf",x"df"),
  1095 => (x"c1",x"80",x"f7",x"50"),
  1096 => (x"c1",x"40",x"e9",x"c3"),
  1097 => (x"ce",x"78",x"f3",x"dd"),
  1098 => (x"cb",x"df",x"c1",x"87"),
  1099 => (x"ec",x"dd",x"c1",x"48"),
  1100 => (x"c1",x"80",x"fc",x"78"),
  1101 => (x"26",x"78",x"c8",x"c4"),
  1102 => (x"5b",x"5e",x"0e",x"4f"),
  1103 => (x"4c",x"71",x"0e",x"5c"),
  1104 => (x"c1",x"92",x"cb",x"4a"),
  1105 => (x"c8",x"82",x"fa",x"dd"),
  1106 => (x"a2",x"c9",x"49",x"a2"),
  1107 => (x"4b",x"6b",x"97",x"4b"),
  1108 => (x"49",x"69",x"97",x"1e"),
  1109 => (x"12",x"82",x"ca",x"1e"),
  1110 => (x"fa",x"e7",x"c0",x"49"),
  1111 => (x"d4",x"49",x"c0",x"87"),
  1112 => (x"49",x"74",x"87",x"c9"),
  1113 => (x"87",x"c1",x"fa",x"c0"),
  1114 => (x"f8",x"f4",x"8e",x"f8"),
  1115 => (x"1e",x"73",x"1e",x"87"),
  1116 => (x"ff",x"49",x"4b",x"71"),
  1117 => (x"49",x"73",x"87",x"c3"),
  1118 => (x"f4",x"87",x"fe",x"fe"),
  1119 => (x"73",x"1e",x"87",x"e9"),
  1120 => (x"c6",x"4b",x"71",x"1e"),
  1121 => (x"db",x"02",x"4a",x"a3"),
  1122 => (x"02",x"8a",x"c1",x"87"),
  1123 => (x"02",x"8a",x"87",x"d6"),
  1124 => (x"8a",x"87",x"da",x"c1"),
  1125 => (x"87",x"fc",x"c0",x"02"),
  1126 => (x"e1",x"c0",x"02",x"8a"),
  1127 => (x"cb",x"02",x"8a",x"87"),
  1128 => (x"87",x"db",x"c1",x"87"),
  1129 => (x"c0",x"fd",x"49",x"c7"),
  1130 => (x"87",x"de",x"c1",x"87"),
  1131 => (x"bf",x"c4",x"ea",x"c2"),
  1132 => (x"87",x"cb",x"c1",x"02"),
  1133 => (x"c2",x"88",x"c1",x"48"),
  1134 => (x"c1",x"58",x"c8",x"ea"),
  1135 => (x"ea",x"c2",x"87",x"c1"),
  1136 => (x"c0",x"02",x"bf",x"c8"),
  1137 => (x"ea",x"c2",x"87",x"f9"),
  1138 => (x"c1",x"48",x"bf",x"c4"),
  1139 => (x"c8",x"ea",x"c2",x"80"),
  1140 => (x"87",x"eb",x"c0",x"58"),
  1141 => (x"bf",x"c4",x"ea",x"c2"),
  1142 => (x"c2",x"89",x"c6",x"49"),
  1143 => (x"c0",x"59",x"c8",x"ea"),
  1144 => (x"da",x"03",x"a9",x"b7"),
  1145 => (x"c4",x"ea",x"c2",x"87"),
  1146 => (x"d2",x"78",x"c0",x"48"),
  1147 => (x"c8",x"ea",x"c2",x"87"),
  1148 => (x"87",x"cb",x"02",x"bf"),
  1149 => (x"bf",x"c4",x"ea",x"c2"),
  1150 => (x"c2",x"80",x"c6",x"48"),
  1151 => (x"c0",x"58",x"c8",x"ea"),
  1152 => (x"87",x"e7",x"d1",x"49"),
  1153 => (x"f7",x"c0",x"49",x"73"),
  1154 => (x"da",x"f2",x"87",x"df"),
  1155 => (x"5b",x"5e",x"0e",x"87"),
  1156 => (x"4c",x"71",x"0e",x"5c"),
  1157 => (x"74",x"1e",x"66",x"cc"),
  1158 => (x"c1",x"93",x"cb",x"4b"),
  1159 => (x"c4",x"83",x"fa",x"dd"),
  1160 => (x"49",x"6a",x"4a",x"a3"),
  1161 => (x"87",x"d0",x"fa",x"fe"),
  1162 => (x"7b",x"e7",x"c2",x"c1"),
  1163 => (x"d4",x"49",x"a3",x"c8"),
  1164 => (x"a3",x"c9",x"51",x"66"),
  1165 => (x"51",x"66",x"d8",x"49"),
  1166 => (x"dc",x"49",x"a3",x"ca"),
  1167 => (x"f1",x"26",x"51",x"66"),
  1168 => (x"5e",x"0e",x"87",x"e3"),
  1169 => (x"0e",x"5d",x"5c",x"5b"),
  1170 => (x"d8",x"86",x"d0",x"ff"),
  1171 => (x"a6",x"c4",x"59",x"a6"),
  1172 => (x"c4",x"78",x"c0",x"48"),
  1173 => (x"66",x"c4",x"c1",x"80"),
  1174 => (x"c1",x"80",x"c4",x"78"),
  1175 => (x"c1",x"80",x"c4",x"78"),
  1176 => (x"c8",x"ea",x"c2",x"78"),
  1177 => (x"c2",x"78",x"c1",x"48"),
  1178 => (x"48",x"bf",x"c0",x"ea"),
  1179 => (x"cb",x"05",x"a8",x"de"),
  1180 => (x"87",x"e5",x"f3",x"87"),
  1181 => (x"a6",x"c8",x"49",x"70"),
  1182 => (x"87",x"f8",x"ce",x"59"),
  1183 => (x"e9",x"87",x"ed",x"e8"),
  1184 => (x"dc",x"e8",x"87",x"cf"),
  1185 => (x"c0",x"4c",x"70",x"87"),
  1186 => (x"c1",x"02",x"ac",x"fb"),
  1187 => (x"66",x"d4",x"87",x"d0"),
  1188 => (x"87",x"c2",x"c1",x"05"),
  1189 => (x"c1",x"1e",x"1e",x"c0"),
  1190 => (x"ed",x"df",x"c1",x"1e"),
  1191 => (x"fd",x"49",x"c0",x"1e"),
  1192 => (x"d0",x"c1",x"87",x"eb"),
  1193 => (x"82",x"c4",x"4a",x"66"),
  1194 => (x"81",x"c7",x"49",x"6a"),
  1195 => (x"1e",x"c1",x"51",x"74"),
  1196 => (x"49",x"6a",x"1e",x"d8"),
  1197 => (x"ec",x"e8",x"81",x"c8"),
  1198 => (x"c1",x"86",x"d8",x"87"),
  1199 => (x"c0",x"48",x"66",x"c4"),
  1200 => (x"87",x"c7",x"01",x"a8"),
  1201 => (x"c1",x"48",x"a6",x"c4"),
  1202 => (x"c1",x"87",x"ce",x"78"),
  1203 => (x"c1",x"48",x"66",x"c4"),
  1204 => (x"58",x"a6",x"cc",x"88"),
  1205 => (x"f8",x"e7",x"87",x"c3"),
  1206 => (x"48",x"a6",x"cc",x"87"),
  1207 => (x"9c",x"74",x"78",x"c2"),
  1208 => (x"87",x"cc",x"cd",x"02"),
  1209 => (x"c1",x"48",x"66",x"c4"),
  1210 => (x"03",x"a8",x"66",x"c8"),
  1211 => (x"d8",x"87",x"c1",x"cd"),
  1212 => (x"78",x"c0",x"48",x"a6"),
  1213 => (x"70",x"87",x"ea",x"e6"),
  1214 => (x"ac",x"d0",x"c1",x"4c"),
  1215 => (x"87",x"d6",x"c2",x"05"),
  1216 => (x"e9",x"7e",x"66",x"d8"),
  1217 => (x"49",x"70",x"87",x"ce"),
  1218 => (x"e6",x"59",x"a6",x"dc"),
  1219 => (x"4c",x"70",x"87",x"d3"),
  1220 => (x"05",x"ac",x"ec",x"c0"),
  1221 => (x"c4",x"87",x"ea",x"c1"),
  1222 => (x"91",x"cb",x"49",x"66"),
  1223 => (x"81",x"66",x"c0",x"c1"),
  1224 => (x"6a",x"4a",x"a1",x"c4"),
  1225 => (x"4a",x"a1",x"c8",x"4d"),
  1226 => (x"c1",x"52",x"66",x"d8"),
  1227 => (x"e5",x"79",x"e9",x"c3"),
  1228 => (x"4c",x"70",x"87",x"ef"),
  1229 => (x"87",x"d8",x"02",x"9c"),
  1230 => (x"02",x"ac",x"fb",x"c0"),
  1231 => (x"55",x"74",x"87",x"d2"),
  1232 => (x"70",x"87",x"de",x"e5"),
  1233 => (x"c7",x"02",x"9c",x"4c"),
  1234 => (x"ac",x"fb",x"c0",x"87"),
  1235 => (x"87",x"ee",x"ff",x"05"),
  1236 => (x"c2",x"55",x"e0",x"c0"),
  1237 => (x"97",x"c0",x"55",x"c1"),
  1238 => (x"49",x"66",x"d4",x"7d"),
  1239 => (x"db",x"05",x"a9",x"6e"),
  1240 => (x"48",x"66",x"c4",x"87"),
  1241 => (x"04",x"a8",x"66",x"c8"),
  1242 => (x"66",x"c4",x"87",x"ca"),
  1243 => (x"c8",x"80",x"c1",x"48"),
  1244 => (x"87",x"c8",x"58",x"a6"),
  1245 => (x"c1",x"48",x"66",x"c8"),
  1246 => (x"58",x"a6",x"cc",x"88"),
  1247 => (x"70",x"87",x"e2",x"e4"),
  1248 => (x"ac",x"d0",x"c1",x"4c"),
  1249 => (x"d0",x"87",x"c8",x"05"),
  1250 => (x"80",x"c1",x"48",x"66"),
  1251 => (x"c1",x"58",x"a6",x"d4"),
  1252 => (x"fd",x"02",x"ac",x"d0"),
  1253 => (x"a6",x"dc",x"87",x"ea"),
  1254 => (x"78",x"66",x"d4",x"48"),
  1255 => (x"dc",x"48",x"66",x"d8"),
  1256 => (x"c9",x"05",x"a8",x"66"),
  1257 => (x"e0",x"c0",x"87",x"dc"),
  1258 => (x"f0",x"c0",x"48",x"a6"),
  1259 => (x"cc",x"80",x"c4",x"78"),
  1260 => (x"80",x"c4",x"78",x"66"),
  1261 => (x"74",x"7e",x"78",x"c0"),
  1262 => (x"88",x"fb",x"c0",x"48"),
  1263 => (x"58",x"a6",x"f0",x"c0"),
  1264 => (x"c8",x"02",x"98",x"70"),
  1265 => (x"cb",x"48",x"87",x"d7"),
  1266 => (x"a6",x"f0",x"c0",x"88"),
  1267 => (x"02",x"98",x"70",x"58"),
  1268 => (x"48",x"87",x"e9",x"c0"),
  1269 => (x"f0",x"c0",x"88",x"c9"),
  1270 => (x"98",x"70",x"58",x"a6"),
  1271 => (x"87",x"e1",x"c3",x"02"),
  1272 => (x"c0",x"88",x"c4",x"48"),
  1273 => (x"70",x"58",x"a6",x"f0"),
  1274 => (x"87",x"de",x"02",x"98"),
  1275 => (x"c0",x"88",x"c1",x"48"),
  1276 => (x"70",x"58",x"a6",x"f0"),
  1277 => (x"c8",x"c3",x"02",x"98"),
  1278 => (x"87",x"db",x"c7",x"87"),
  1279 => (x"48",x"a6",x"e0",x"c0"),
  1280 => (x"66",x"cc",x"78",x"c0"),
  1281 => (x"d0",x"80",x"c1",x"48"),
  1282 => (x"d4",x"e2",x"58",x"a6"),
  1283 => (x"c0",x"4c",x"70",x"87"),
  1284 => (x"d5",x"02",x"ac",x"ec"),
  1285 => (x"66",x"e0",x"c0",x"87"),
  1286 => (x"c0",x"87",x"c6",x"02"),
  1287 => (x"c9",x"5c",x"a6",x"e4"),
  1288 => (x"c0",x"48",x"74",x"87"),
  1289 => (x"e8",x"c0",x"88",x"f0"),
  1290 => (x"ec",x"c0",x"58",x"a6"),
  1291 => (x"87",x"cc",x"02",x"ac"),
  1292 => (x"70",x"87",x"ee",x"e1"),
  1293 => (x"ac",x"ec",x"c0",x"4c"),
  1294 => (x"87",x"f4",x"ff",x"05"),
  1295 => (x"1e",x"66",x"e0",x"c0"),
  1296 => (x"1e",x"49",x"66",x"d4"),
  1297 => (x"1e",x"66",x"ec",x"c0"),
  1298 => (x"1e",x"ed",x"df",x"c1"),
  1299 => (x"f6",x"49",x"66",x"d4"),
  1300 => (x"1e",x"c0",x"87",x"fb"),
  1301 => (x"66",x"dc",x"1e",x"ca"),
  1302 => (x"c1",x"91",x"cb",x"49"),
  1303 => (x"d8",x"81",x"66",x"d8"),
  1304 => (x"a1",x"c4",x"48",x"a6"),
  1305 => (x"bf",x"66",x"d8",x"78"),
  1306 => (x"87",x"f9",x"e1",x"49"),
  1307 => (x"b7",x"c0",x"86",x"d8"),
  1308 => (x"c7",x"c1",x"06",x"a8"),
  1309 => (x"de",x"1e",x"c1",x"87"),
  1310 => (x"bf",x"66",x"c8",x"1e"),
  1311 => (x"87",x"e5",x"e1",x"49"),
  1312 => (x"49",x"70",x"86",x"c8"),
  1313 => (x"88",x"08",x"c0",x"48"),
  1314 => (x"58",x"a6",x"e4",x"c0"),
  1315 => (x"06",x"a8",x"b7",x"c0"),
  1316 => (x"c0",x"87",x"e9",x"c0"),
  1317 => (x"dd",x"48",x"66",x"e0"),
  1318 => (x"df",x"03",x"a8",x"b7"),
  1319 => (x"49",x"bf",x"6e",x"87"),
  1320 => (x"81",x"66",x"e0",x"c0"),
  1321 => (x"66",x"51",x"e0",x"c0"),
  1322 => (x"6e",x"81",x"c1",x"49"),
  1323 => (x"c1",x"c2",x"81",x"bf"),
  1324 => (x"66",x"e0",x"c0",x"51"),
  1325 => (x"6e",x"81",x"c2",x"49"),
  1326 => (x"51",x"c0",x"81",x"bf"),
  1327 => (x"dc",x"c4",x"7e",x"c1"),
  1328 => (x"87",x"d0",x"e2",x"87"),
  1329 => (x"58",x"a6",x"e4",x"c0"),
  1330 => (x"c0",x"87",x"c9",x"e2"),
  1331 => (x"c0",x"58",x"a6",x"e8"),
  1332 => (x"c0",x"05",x"a8",x"ec"),
  1333 => (x"e4",x"c0",x"87",x"cb"),
  1334 => (x"e0",x"c0",x"48",x"a6"),
  1335 => (x"c4",x"c0",x"78",x"66"),
  1336 => (x"fc",x"de",x"ff",x"87"),
  1337 => (x"49",x"66",x"c4",x"87"),
  1338 => (x"c0",x"c1",x"91",x"cb"),
  1339 => (x"80",x"71",x"48",x"66"),
  1340 => (x"4a",x"6e",x"7e",x"70"),
  1341 => (x"49",x"6e",x"82",x"c8"),
  1342 => (x"e0",x"c0",x"81",x"ca"),
  1343 => (x"e4",x"c0",x"51",x"66"),
  1344 => (x"81",x"c1",x"49",x"66"),
  1345 => (x"89",x"66",x"e0",x"c0"),
  1346 => (x"30",x"71",x"48",x"c1"),
  1347 => (x"89",x"c1",x"49",x"70"),
  1348 => (x"c2",x"7a",x"97",x"71"),
  1349 => (x"49",x"bf",x"f5",x"ed"),
  1350 => (x"29",x"66",x"e0",x"c0"),
  1351 => (x"48",x"4a",x"6a",x"97"),
  1352 => (x"f0",x"c0",x"98",x"71"),
  1353 => (x"49",x"6e",x"58",x"a6"),
  1354 => (x"4d",x"69",x"81",x"c4"),
  1355 => (x"d8",x"48",x"66",x"dc"),
  1356 => (x"c0",x"02",x"a8",x"66"),
  1357 => (x"a6",x"d8",x"87",x"c8"),
  1358 => (x"c0",x"78",x"c0",x"48"),
  1359 => (x"a6",x"d8",x"87",x"c5"),
  1360 => (x"d8",x"78",x"c1",x"48"),
  1361 => (x"e0",x"c0",x"1e",x"66"),
  1362 => (x"ff",x"49",x"75",x"1e"),
  1363 => (x"c8",x"87",x"d6",x"de"),
  1364 => (x"c0",x"4c",x"70",x"86"),
  1365 => (x"c1",x"06",x"ac",x"b7"),
  1366 => (x"85",x"74",x"87",x"d4"),
  1367 => (x"74",x"49",x"e0",x"c0"),
  1368 => (x"c1",x"4b",x"75",x"89"),
  1369 => (x"71",x"4a",x"e8",x"d9"),
  1370 => (x"87",x"fc",x"ec",x"fe"),
  1371 => (x"e8",x"c0",x"85",x"c2"),
  1372 => (x"80",x"c1",x"48",x"66"),
  1373 => (x"58",x"a6",x"ec",x"c0"),
  1374 => (x"49",x"66",x"ec",x"c0"),
  1375 => (x"a9",x"70",x"81",x"c1"),
  1376 => (x"87",x"c8",x"c0",x"02"),
  1377 => (x"c0",x"48",x"a6",x"d8"),
  1378 => (x"87",x"c5",x"c0",x"78"),
  1379 => (x"c1",x"48",x"a6",x"d8"),
  1380 => (x"1e",x"66",x"d8",x"78"),
  1381 => (x"c0",x"49",x"a4",x"c2"),
  1382 => (x"88",x"71",x"48",x"e0"),
  1383 => (x"75",x"1e",x"49",x"70"),
  1384 => (x"c0",x"dd",x"ff",x"49"),
  1385 => (x"c0",x"86",x"c8",x"87"),
  1386 => (x"ff",x"01",x"a8",x"b7"),
  1387 => (x"e8",x"c0",x"87",x"c0"),
  1388 => (x"d1",x"c0",x"02",x"66"),
  1389 => (x"c9",x"49",x"6e",x"87"),
  1390 => (x"66",x"e8",x"c0",x"81"),
  1391 => (x"c1",x"48",x"6e",x"51"),
  1392 => (x"c0",x"78",x"f9",x"c4"),
  1393 => (x"49",x"6e",x"87",x"cc"),
  1394 => (x"51",x"c2",x"81",x"c9"),
  1395 => (x"c5",x"c1",x"48",x"6e"),
  1396 => (x"7e",x"c1",x"78",x"ed"),
  1397 => (x"ff",x"87",x"c6",x"c0"),
  1398 => (x"70",x"87",x"f6",x"db"),
  1399 => (x"c0",x"02",x"6e",x"4c"),
  1400 => (x"66",x"c4",x"87",x"f5"),
  1401 => (x"a8",x"66",x"c8",x"48"),
  1402 => (x"87",x"cb",x"c0",x"04"),
  1403 => (x"c1",x"48",x"66",x"c4"),
  1404 => (x"58",x"a6",x"c8",x"80"),
  1405 => (x"c8",x"87",x"e0",x"c0"),
  1406 => (x"88",x"c1",x"48",x"66"),
  1407 => (x"c0",x"58",x"a6",x"cc"),
  1408 => (x"c6",x"c1",x"87",x"d5"),
  1409 => (x"c8",x"c0",x"05",x"ac"),
  1410 => (x"48",x"66",x"cc",x"87"),
  1411 => (x"a6",x"d0",x"80",x"c1"),
  1412 => (x"fc",x"da",x"ff",x"58"),
  1413 => (x"d0",x"4c",x"70",x"87"),
  1414 => (x"80",x"c1",x"48",x"66"),
  1415 => (x"74",x"58",x"a6",x"d4"),
  1416 => (x"cb",x"c0",x"02",x"9c"),
  1417 => (x"48",x"66",x"c4",x"87"),
  1418 => (x"a8",x"66",x"c8",x"c1"),
  1419 => (x"87",x"ff",x"f2",x"04"),
  1420 => (x"87",x"d4",x"da",x"ff"),
  1421 => (x"c7",x"48",x"66",x"c4"),
  1422 => (x"e5",x"c0",x"03",x"a8"),
  1423 => (x"c8",x"ea",x"c2",x"87"),
  1424 => (x"c4",x"78",x"c0",x"48"),
  1425 => (x"91",x"cb",x"49",x"66"),
  1426 => (x"81",x"66",x"c0",x"c1"),
  1427 => (x"6a",x"4a",x"a1",x"c4"),
  1428 => (x"79",x"52",x"c0",x"4a"),
  1429 => (x"c1",x"48",x"66",x"c4"),
  1430 => (x"58",x"a6",x"c8",x"80"),
  1431 => (x"ff",x"04",x"a8",x"c7"),
  1432 => (x"d0",x"ff",x"87",x"db"),
  1433 => (x"87",x"fb",x"e0",x"8e"),
  1434 => (x"1e",x"00",x"20",x"3a"),
  1435 => (x"4b",x"71",x"1e",x"73"),
  1436 => (x"87",x"c6",x"02",x"9b"),
  1437 => (x"48",x"c4",x"ea",x"c2"),
  1438 => (x"1e",x"c7",x"78",x"c0"),
  1439 => (x"bf",x"c4",x"ea",x"c2"),
  1440 => (x"dd",x"c1",x"1e",x"49"),
  1441 => (x"ea",x"c2",x"1e",x"fa"),
  1442 => (x"ee",x"49",x"bf",x"c0"),
  1443 => (x"86",x"cc",x"87",x"f4"),
  1444 => (x"bf",x"c0",x"ea",x"c2"),
  1445 => (x"87",x"f9",x"e9",x"49"),
  1446 => (x"c8",x"02",x"9b",x"73"),
  1447 => (x"fa",x"dd",x"c1",x"87"),
  1448 => (x"d6",x"e6",x"c0",x"49"),
  1449 => (x"fe",x"df",x"ff",x"87"),
  1450 => (x"1e",x"73",x"1e",x"87"),
  1451 => (x"db",x"c2",x"4b",x"c0"),
  1452 => (x"50",x"c0",x"48",x"d2"),
  1453 => (x"bf",x"dd",x"df",x"c1"),
  1454 => (x"ea",x"fb",x"c0",x"49"),
  1455 => (x"05",x"98",x"70",x"87"),
  1456 => (x"db",x"c1",x"87",x"c4"),
  1457 => (x"48",x"73",x"4b",x"cc"),
  1458 => (x"87",x"db",x"df",x"ff"),
  1459 => (x"20",x"4d",x"4f",x"52"),
  1460 => (x"64",x"61",x"6f",x"6c"),
  1461 => (x"20",x"67",x"6e",x"69"),
  1462 => (x"6c",x"69",x"61",x"66"),
  1463 => (x"1e",x"00",x"64",x"65"),
  1464 => (x"c1",x"87",x"e9",x"c7"),
  1465 => (x"87",x"c3",x"fe",x"49"),
  1466 => (x"87",x"cf",x"ef",x"fe"),
  1467 => (x"cd",x"02",x"98",x"70"),
  1468 => (x"cc",x"f8",x"fe",x"87"),
  1469 => (x"02",x"98",x"70",x"87"),
  1470 => (x"4a",x"c1",x"87",x"c4"),
  1471 => (x"4a",x"c0",x"87",x"c2"),
  1472 => (x"ce",x"05",x"9a",x"72"),
  1473 => (x"c1",x"1e",x"c0",x"87"),
  1474 => (x"c0",x"49",x"f3",x"dc"),
  1475 => (x"c4",x"87",x"fb",x"f0"),
  1476 => (x"c0",x"87",x"fe",x"86"),
  1477 => (x"c0",x"87",x"e5",x"ff"),
  1478 => (x"fe",x"dc",x"c1",x"1e"),
  1479 => (x"e9",x"f0",x"c0",x"49"),
  1480 => (x"fe",x"1e",x"c0",x"87"),
  1481 => (x"49",x"70",x"87",x"c3"),
  1482 => (x"87",x"de",x"f0",x"c0"),
  1483 => (x"f8",x"87",x"dc",x"c3"),
  1484 => (x"53",x"4f",x"26",x"8e"),
  1485 => (x"61",x"66",x"20",x"44"),
  1486 => (x"64",x"65",x"6c",x"69"),
  1487 => (x"6f",x"42",x"00",x"2e"),
  1488 => (x"6e",x"69",x"74",x"6f"),
  1489 => (x"2e",x"2e",x"2e",x"67"),
  1490 => (x"e8",x"c0",x"1e",x"00"),
  1491 => (x"f3",x"c0",x"87",x"c9"),
  1492 => (x"87",x"f6",x"87",x"ee"),
  1493 => (x"c2",x"1e",x"4f",x"26"),
  1494 => (x"c0",x"48",x"c4",x"ea"),
  1495 => (x"c0",x"ea",x"c2",x"78"),
  1496 => (x"fd",x"78",x"c0",x"48"),
  1497 => (x"87",x"e1",x"87",x"f9"),
  1498 => (x"4f",x"26",x"48",x"c0"),
  1499 => (x"78",x"45",x"20",x"80"),
  1500 => (x"80",x"00",x"74",x"69"),
  1501 => (x"63",x"61",x"42",x"20"),
  1502 => (x"10",x"e9",x"00",x"6b"),
  1503 => (x"2a",x"99",x"00",x"00"),
  1504 => (x"00",x"00",x"00",x"00"),
  1505 => (x"00",x"10",x"e9",x"00"),
  1506 => (x"00",x"2a",x"b7",x"00"),
  1507 => (x"00",x"00",x"00",x"00"),
  1508 => (x"00",x"00",x"10",x"e9"),
  1509 => (x"00",x"00",x"2a",x"d5"),
  1510 => (x"e9",x"00",x"00",x"00"),
  1511 => (x"f3",x"00",x"00",x"10"),
  1512 => (x"00",x"00",x"00",x"2a"),
  1513 => (x"10",x"e9",x"00",x"00"),
  1514 => (x"2b",x"11",x"00",x"00"),
  1515 => (x"00",x"00",x"00",x"00"),
  1516 => (x"00",x"10",x"e9",x"00"),
  1517 => (x"00",x"2b",x"2f",x"00"),
  1518 => (x"00",x"00",x"00",x"00"),
  1519 => (x"00",x"00",x"10",x"e9"),
  1520 => (x"00",x"00",x"2b",x"4d"),
  1521 => (x"e9",x"00",x"00",x"00"),
  1522 => (x"00",x"00",x"00",x"10"),
  1523 => (x"00",x"00",x"00",x"00"),
  1524 => (x"11",x"7e",x"00",x"00"),
  1525 => (x"00",x"00",x"00",x"00"),
  1526 => (x"00",x"00",x"00",x"00"),
  1527 => (x"00",x"17",x"e1",x"00"),
  1528 => (x"53",x"4d",x"41",x"00"),
  1529 => (x"44",x"41",x"52",x"54"),
  1530 => (x"4d",x"4f",x"52",x"20"),
  1531 => (x"61",x"6f",x"4c",x"00"),
  1532 => (x"2e",x"2a",x"20",x"64"),
  1533 => (x"f0",x"fe",x"1e",x"00"),
  1534 => (x"cd",x"78",x"c0",x"48"),
  1535 => (x"26",x"09",x"79",x"09"),
  1536 => (x"fe",x"1e",x"1e",x"4f"),
  1537 => (x"48",x"7e",x"bf",x"f0"),
  1538 => (x"1e",x"4f",x"26",x"26"),
  1539 => (x"c1",x"48",x"f0",x"fe"),
  1540 => (x"1e",x"4f",x"26",x"78"),
  1541 => (x"c0",x"48",x"f0",x"fe"),
  1542 => (x"1e",x"4f",x"26",x"78"),
  1543 => (x"52",x"c0",x"4a",x"71"),
  1544 => (x"0e",x"4f",x"26",x"52"),
  1545 => (x"5d",x"5c",x"5b",x"5e"),
  1546 => (x"71",x"86",x"f4",x"0e"),
  1547 => (x"7e",x"6d",x"97",x"4d"),
  1548 => (x"97",x"4c",x"a5",x"c1"),
  1549 => (x"a6",x"c8",x"48",x"6c"),
  1550 => (x"c4",x"48",x"6e",x"58"),
  1551 => (x"c5",x"05",x"a8",x"66"),
  1552 => (x"c0",x"48",x"ff",x"87"),
  1553 => (x"ca",x"ff",x"87",x"e6"),
  1554 => (x"49",x"a5",x"c2",x"87"),
  1555 => (x"71",x"4b",x"6c",x"97"),
  1556 => (x"6b",x"97",x"4b",x"a3"),
  1557 => (x"7e",x"6c",x"97",x"4b"),
  1558 => (x"80",x"c1",x"48",x"6e"),
  1559 => (x"c7",x"58",x"a6",x"c8"),
  1560 => (x"58",x"a6",x"cc",x"98"),
  1561 => (x"fe",x"7c",x"97",x"70"),
  1562 => (x"48",x"73",x"87",x"e1"),
  1563 => (x"4d",x"26",x"8e",x"f4"),
  1564 => (x"4b",x"26",x"4c",x"26"),
  1565 => (x"5e",x"0e",x"4f",x"26"),
  1566 => (x"f4",x"0e",x"5c",x"5b"),
  1567 => (x"d8",x"4c",x"71",x"86"),
  1568 => (x"ff",x"c3",x"4a",x"66"),
  1569 => (x"4b",x"a4",x"c2",x"9a"),
  1570 => (x"73",x"49",x"6c",x"97"),
  1571 => (x"51",x"72",x"49",x"a1"),
  1572 => (x"6e",x"7e",x"6c",x"97"),
  1573 => (x"c8",x"80",x"c1",x"48"),
  1574 => (x"98",x"c7",x"58",x"a6"),
  1575 => (x"70",x"58",x"a6",x"cc"),
  1576 => (x"ff",x"8e",x"f4",x"54"),
  1577 => (x"1e",x"1e",x"87",x"ca"),
  1578 => (x"e0",x"87",x"e8",x"fd"),
  1579 => (x"c0",x"49",x"4a",x"bf"),
  1580 => (x"02",x"99",x"c0",x"e0"),
  1581 => (x"1e",x"72",x"87",x"cb"),
  1582 => (x"49",x"eb",x"ed",x"c2"),
  1583 => (x"c4",x"87",x"f7",x"fe"),
  1584 => (x"87",x"fd",x"fc",x"86"),
  1585 => (x"c2",x"fd",x"7e",x"70"),
  1586 => (x"4f",x"26",x"26",x"87"),
  1587 => (x"eb",x"ed",x"c2",x"1e"),
  1588 => (x"87",x"c7",x"fd",x"49"),
  1589 => (x"49",x"e6",x"e2",x"c1"),
  1590 => (x"c5",x"87",x"da",x"fc"),
  1591 => (x"4f",x"26",x"87",x"d9"),
  1592 => (x"5c",x"5b",x"5e",x"0e"),
  1593 => (x"ee",x"c2",x"0e",x"5d"),
  1594 => (x"c1",x"4a",x"bf",x"ca"),
  1595 => (x"49",x"bf",x"f4",x"e4"),
  1596 => (x"71",x"bc",x"72",x"4c"),
  1597 => (x"87",x"db",x"fc",x"4d"),
  1598 => (x"49",x"74",x"4b",x"c0"),
  1599 => (x"d5",x"02",x"99",x"d0"),
  1600 => (x"d0",x"49",x"75",x"87"),
  1601 => (x"c0",x"1e",x"71",x"99"),
  1602 => (x"c6",x"eb",x"c1",x"1e"),
  1603 => (x"12",x"82",x"73",x"4a"),
  1604 => (x"87",x"e4",x"c0",x"49"),
  1605 => (x"2c",x"c1",x"86",x"c8"),
  1606 => (x"ab",x"c8",x"83",x"2d"),
  1607 => (x"87",x"da",x"ff",x"04"),
  1608 => (x"c1",x"87",x"e8",x"fb"),
  1609 => (x"c2",x"48",x"f4",x"e4"),
  1610 => (x"78",x"bf",x"ca",x"ee"),
  1611 => (x"4c",x"26",x"4d",x"26"),
  1612 => (x"4f",x"26",x"4b",x"26"),
  1613 => (x"00",x"00",x"00",x"00"),
  1614 => (x"48",x"d0",x"ff",x"1e"),
  1615 => (x"ff",x"78",x"e1",x"c8"),
  1616 => (x"78",x"c5",x"48",x"d4"),
  1617 => (x"c3",x"02",x"66",x"c4"),
  1618 => (x"78",x"e0",x"c3",x"87"),
  1619 => (x"c6",x"02",x"66",x"c8"),
  1620 => (x"48",x"d4",x"ff",x"87"),
  1621 => (x"ff",x"78",x"f0",x"c3"),
  1622 => (x"78",x"71",x"48",x"d4"),
  1623 => (x"c8",x"48",x"d0",x"ff"),
  1624 => (x"e0",x"c0",x"78",x"e1"),
  1625 => (x"0e",x"4f",x"26",x"78"),
  1626 => (x"0e",x"5c",x"5b",x"5e"),
  1627 => (x"ed",x"c2",x"4c",x"71"),
  1628 => (x"ee",x"fa",x"49",x"eb"),
  1629 => (x"c0",x"4a",x"70",x"87"),
  1630 => (x"c2",x"04",x"aa",x"b7"),
  1631 => (x"e0",x"c3",x"87",x"e3"),
  1632 => (x"87",x"c9",x"05",x"aa"),
  1633 => (x"48",x"ea",x"e8",x"c1"),
  1634 => (x"d4",x"c2",x"78",x"c1"),
  1635 => (x"aa",x"f0",x"c3",x"87"),
  1636 => (x"c1",x"87",x"c9",x"05"),
  1637 => (x"c1",x"48",x"e6",x"e8"),
  1638 => (x"87",x"f5",x"c1",x"78"),
  1639 => (x"bf",x"ea",x"e8",x"c1"),
  1640 => (x"72",x"87",x"c7",x"02"),
  1641 => (x"b3",x"c0",x"c2",x"4b"),
  1642 => (x"4b",x"72",x"87",x"c2"),
  1643 => (x"d1",x"05",x"9c",x"74"),
  1644 => (x"e6",x"e8",x"c1",x"87"),
  1645 => (x"e8",x"c1",x"1e",x"bf"),
  1646 => (x"72",x"1e",x"bf",x"ea"),
  1647 => (x"87",x"f8",x"fd",x"49"),
  1648 => (x"e8",x"c1",x"86",x"c8"),
  1649 => (x"c0",x"02",x"bf",x"e6"),
  1650 => (x"49",x"73",x"87",x"e0"),
  1651 => (x"91",x"29",x"b7",x"c4"),
  1652 => (x"81",x"c6",x"ea",x"c1"),
  1653 => (x"9a",x"cf",x"4a",x"73"),
  1654 => (x"48",x"c1",x"92",x"c2"),
  1655 => (x"4a",x"70",x"30",x"72"),
  1656 => (x"48",x"72",x"ba",x"ff"),
  1657 => (x"79",x"70",x"98",x"69"),
  1658 => (x"49",x"73",x"87",x"db"),
  1659 => (x"91",x"29",x"b7",x"c4"),
  1660 => (x"81",x"c6",x"ea",x"c1"),
  1661 => (x"9a",x"cf",x"4a",x"73"),
  1662 => (x"48",x"c3",x"92",x"c2"),
  1663 => (x"4a",x"70",x"30",x"72"),
  1664 => (x"70",x"b0",x"69",x"48"),
  1665 => (x"ea",x"e8",x"c1",x"79"),
  1666 => (x"c1",x"78",x"c0",x"48"),
  1667 => (x"c0",x"48",x"e6",x"e8"),
  1668 => (x"eb",x"ed",x"c2",x"78"),
  1669 => (x"87",x"cb",x"f8",x"49"),
  1670 => (x"b7",x"c0",x"4a",x"70"),
  1671 => (x"dd",x"fd",x"03",x"aa"),
  1672 => (x"fc",x"48",x"c0",x"87"),
  1673 => (x"00",x"00",x"87",x"c8"),
  1674 => (x"00",x"00",x"00",x"00"),
  1675 => (x"71",x"1e",x"00",x"00"),
  1676 => (x"f2",x"fc",x"49",x"4a"),
  1677 => (x"1e",x"4f",x"26",x"87"),
  1678 => (x"49",x"72",x"4a",x"c0"),
  1679 => (x"ea",x"c1",x"91",x"c4"),
  1680 => (x"79",x"c0",x"81",x"c6"),
  1681 => (x"b7",x"d0",x"82",x"c1"),
  1682 => (x"87",x"ee",x"04",x"aa"),
  1683 => (x"5e",x"0e",x"4f",x"26"),
  1684 => (x"0e",x"5d",x"5c",x"5b"),
  1685 => (x"fa",x"f6",x"4d",x"71"),
  1686 => (x"c4",x"4a",x"75",x"87"),
  1687 => (x"c1",x"92",x"2a",x"b7"),
  1688 => (x"75",x"82",x"c6",x"ea"),
  1689 => (x"c2",x"9c",x"cf",x"4c"),
  1690 => (x"4b",x"49",x"6a",x"94"),
  1691 => (x"9b",x"c3",x"2b",x"74"),
  1692 => (x"30",x"74",x"48",x"c2"),
  1693 => (x"bc",x"ff",x"4c",x"70"),
  1694 => (x"98",x"71",x"48",x"74"),
  1695 => (x"ca",x"f6",x"7a",x"70"),
  1696 => (x"fa",x"48",x"73",x"87"),
  1697 => (x"00",x"00",x"87",x"e6"),
  1698 => (x"00",x"00",x"00",x"00"),
  1699 => (x"00",x"00",x"00",x"00"),
  1700 => (x"00",x"00",x"00",x"00"),
  1701 => (x"00",x"00",x"00",x"00"),
  1702 => (x"00",x"00",x"00",x"00"),
  1703 => (x"00",x"00",x"00",x"00"),
  1704 => (x"00",x"00",x"00",x"00"),
  1705 => (x"00",x"00",x"00",x"00"),
  1706 => (x"00",x"00",x"00",x"00"),
  1707 => (x"00",x"00",x"00",x"00"),
  1708 => (x"00",x"00",x"00",x"00"),
  1709 => (x"00",x"00",x"00",x"00"),
  1710 => (x"00",x"00",x"00",x"00"),
  1711 => (x"00",x"00",x"00",x"00"),
  1712 => (x"00",x"00",x"00",x"00"),
  1713 => (x"1e",x"16",x"00",x"00"),
  1714 => (x"36",x"2e",x"25",x"26"),
  1715 => (x"ff",x"1e",x"3e",x"3d"),
  1716 => (x"e1",x"c8",x"48",x"d0"),
  1717 => (x"ff",x"48",x"71",x"78"),
  1718 => (x"26",x"78",x"08",x"d4"),
  1719 => (x"d0",x"ff",x"1e",x"4f"),
  1720 => (x"78",x"e1",x"c8",x"48"),
  1721 => (x"d4",x"ff",x"48",x"71"),
  1722 => (x"66",x"c4",x"78",x"08"),
  1723 => (x"08",x"d4",x"ff",x"48"),
  1724 => (x"1e",x"4f",x"26",x"78"),
  1725 => (x"66",x"c4",x"4a",x"71"),
  1726 => (x"49",x"72",x"1e",x"49"),
  1727 => (x"ff",x"87",x"de",x"ff"),
  1728 => (x"e0",x"c0",x"48",x"d0"),
  1729 => (x"4f",x"26",x"26",x"78"),
  1730 => (x"c4",x"4a",x"71",x"1e"),
  1731 => (x"e0",x"c1",x"1e",x"66"),
  1732 => (x"c8",x"ff",x"49",x"a2"),
  1733 => (x"49",x"66",x"c8",x"87"),
  1734 => (x"ff",x"29",x"b7",x"c8"),
  1735 => (x"78",x"71",x"48",x"d4"),
  1736 => (x"c0",x"48",x"d0",x"ff"),
  1737 => (x"26",x"26",x"78",x"e0"),
  1738 => (x"d4",x"ff",x"1e",x"4f"),
  1739 => (x"7a",x"ff",x"c3",x"4a"),
  1740 => (x"c8",x"48",x"d0",x"ff"),
  1741 => (x"7a",x"de",x"78",x"e1"),
  1742 => (x"bf",x"f5",x"ed",x"c2"),
  1743 => (x"c8",x"48",x"49",x"7a"),
  1744 => (x"71",x"7a",x"70",x"28"),
  1745 => (x"70",x"28",x"d0",x"48"),
  1746 => (x"d8",x"48",x"71",x"7a"),
  1747 => (x"ff",x"7a",x"70",x"28"),
  1748 => (x"e0",x"c0",x"48",x"d0"),
  1749 => (x"0e",x"4f",x"26",x"78"),
  1750 => (x"5d",x"5c",x"5b",x"5e"),
  1751 => (x"c2",x"4c",x"71",x"0e"),
  1752 => (x"4d",x"bf",x"f5",x"ed"),
  1753 => (x"d0",x"2b",x"74",x"4b"),
  1754 => (x"83",x"c1",x"9b",x"66"),
  1755 => (x"04",x"ab",x"66",x"d4"),
  1756 => (x"4b",x"c0",x"87",x"c2"),
  1757 => (x"66",x"d0",x"4a",x"74"),
  1758 => (x"ff",x"31",x"72",x"49"),
  1759 => (x"73",x"99",x"75",x"b9"),
  1760 => (x"70",x"30",x"72",x"48"),
  1761 => (x"b0",x"71",x"48",x"4a"),
  1762 => (x"58",x"f9",x"ed",x"c2"),
  1763 => (x"26",x"87",x"da",x"fe"),
  1764 => (x"26",x"4c",x"26",x"4d"),
  1765 => (x"1e",x"4f",x"26",x"4b"),
  1766 => (x"c8",x"48",x"d0",x"ff"),
  1767 => (x"48",x"71",x"78",x"c9"),
  1768 => (x"78",x"08",x"d4",x"ff"),
  1769 => (x"71",x"1e",x"4f",x"26"),
  1770 => (x"87",x"eb",x"49",x"4a"),
  1771 => (x"c8",x"48",x"d0",x"ff"),
  1772 => (x"1e",x"4f",x"26",x"78"),
  1773 => (x"4b",x"71",x"1e",x"73"),
  1774 => (x"bf",x"c5",x"ee",x"c2"),
  1775 => (x"c2",x"87",x"c3",x"02"),
  1776 => (x"d0",x"ff",x"87",x"eb"),
  1777 => (x"78",x"c9",x"c8",x"48"),
  1778 => (x"e0",x"c0",x"49",x"73"),
  1779 => (x"48",x"d4",x"ff",x"b1"),
  1780 => (x"ed",x"c2",x"78",x"71"),
  1781 => (x"78",x"c0",x"48",x"f9"),
  1782 => (x"c5",x"02",x"66",x"c8"),
  1783 => (x"49",x"ff",x"c3",x"87"),
  1784 => (x"49",x"c0",x"87",x"c2"),
  1785 => (x"59",x"c1",x"ee",x"c2"),
  1786 => (x"c6",x"02",x"66",x"cc"),
  1787 => (x"d5",x"d5",x"c5",x"87"),
  1788 => (x"cf",x"87",x"c4",x"4a"),
  1789 => (x"c2",x"4a",x"ff",x"ff"),
  1790 => (x"c2",x"5a",x"c5",x"ee"),
  1791 => (x"c1",x"48",x"c5",x"ee"),
  1792 => (x"26",x"87",x"c4",x"78"),
  1793 => (x"26",x"4c",x"26",x"4d"),
  1794 => (x"0e",x"4f",x"26",x"4b"),
  1795 => (x"5d",x"5c",x"5b",x"5e"),
  1796 => (x"c2",x"4a",x"71",x"0e"),
  1797 => (x"4c",x"bf",x"c1",x"ee"),
  1798 => (x"cb",x"02",x"9a",x"72"),
  1799 => (x"91",x"c8",x"49",x"87"),
  1800 => (x"4b",x"e9",x"ee",x"c1"),
  1801 => (x"87",x"c4",x"83",x"71"),
  1802 => (x"4b",x"e9",x"f2",x"c1"),
  1803 => (x"49",x"13",x"4d",x"c0"),
  1804 => (x"ed",x"c2",x"99",x"74"),
  1805 => (x"ff",x"b9",x"bf",x"fd"),
  1806 => (x"78",x"71",x"48",x"d4"),
  1807 => (x"85",x"2c",x"b7",x"c1"),
  1808 => (x"04",x"ad",x"b7",x"c8"),
  1809 => (x"ed",x"c2",x"87",x"e8"),
  1810 => (x"c8",x"48",x"bf",x"f9"),
  1811 => (x"fd",x"ed",x"c2",x"80"),
  1812 => (x"87",x"ef",x"fe",x"58"),
  1813 => (x"71",x"1e",x"73",x"1e"),
  1814 => (x"9a",x"4a",x"13",x"4b"),
  1815 => (x"72",x"87",x"cb",x"02"),
  1816 => (x"87",x"e7",x"fe",x"49"),
  1817 => (x"05",x"9a",x"4a",x"13"),
  1818 => (x"da",x"fe",x"87",x"f5"),
  1819 => (x"ed",x"c2",x"1e",x"87"),
  1820 => (x"c2",x"49",x"bf",x"f9"),
  1821 => (x"c1",x"48",x"f9",x"ed"),
  1822 => (x"c0",x"c4",x"78",x"a1"),
  1823 => (x"db",x"03",x"a9",x"b7"),
  1824 => (x"48",x"d4",x"ff",x"87"),
  1825 => (x"bf",x"fd",x"ed",x"c2"),
  1826 => (x"f9",x"ed",x"c2",x"78"),
  1827 => (x"ed",x"c2",x"49",x"bf"),
  1828 => (x"a1",x"c1",x"48",x"f9"),
  1829 => (x"b7",x"c0",x"c4",x"78"),
  1830 => (x"87",x"e5",x"04",x"a9"),
  1831 => (x"c8",x"48",x"d0",x"ff"),
  1832 => (x"c5",x"ee",x"c2",x"78"),
  1833 => (x"26",x"78",x"c0",x"48"),
  1834 => (x"00",x"00",x"00",x"4f"),
  1835 => (x"00",x"00",x"00",x"00"),
  1836 => (x"00",x"00",x"00",x"00"),
  1837 => (x"00",x"00",x"5f",x"5f"),
  1838 => (x"03",x"03",x"00",x"00"),
  1839 => (x"00",x"03",x"03",x"00"),
  1840 => (x"7f",x"7f",x"14",x"00"),
  1841 => (x"14",x"7f",x"7f",x"14"),
  1842 => (x"2e",x"24",x"00",x"00"),
  1843 => (x"12",x"3a",x"6b",x"6b"),
  1844 => (x"36",x"6a",x"4c",x"00"),
  1845 => (x"32",x"56",x"6c",x"18"),
  1846 => (x"4f",x"7e",x"30",x"00"),
  1847 => (x"68",x"3a",x"77",x"59"),
  1848 => (x"04",x"00",x"00",x"40"),
  1849 => (x"00",x"00",x"03",x"07"),
  1850 => (x"1c",x"00",x"00",x"00"),
  1851 => (x"00",x"41",x"63",x"3e"),
  1852 => (x"41",x"00",x"00",x"00"),
  1853 => (x"00",x"1c",x"3e",x"63"),
  1854 => (x"3e",x"2a",x"08",x"00"),
  1855 => (x"2a",x"3e",x"1c",x"1c"),
  1856 => (x"08",x"08",x"00",x"08"),
  1857 => (x"08",x"08",x"3e",x"3e"),
  1858 => (x"80",x"00",x"00",x"00"),
  1859 => (x"00",x"00",x"60",x"e0"),
  1860 => (x"08",x"08",x"00",x"00"),
  1861 => (x"08",x"08",x"08",x"08"),
  1862 => (x"00",x"00",x"00",x"00"),
  1863 => (x"00",x"00",x"60",x"60"),
  1864 => (x"30",x"60",x"40",x"00"),
  1865 => (x"03",x"06",x"0c",x"18"),
  1866 => (x"7f",x"3e",x"00",x"01"),
  1867 => (x"3e",x"7f",x"4d",x"59"),
  1868 => (x"06",x"04",x"00",x"00"),
  1869 => (x"00",x"00",x"7f",x"7f"),
  1870 => (x"63",x"42",x"00",x"00"),
  1871 => (x"46",x"4f",x"59",x"71"),
  1872 => (x"63",x"22",x"00",x"00"),
  1873 => (x"36",x"7f",x"49",x"49"),
  1874 => (x"16",x"1c",x"18",x"00"),
  1875 => (x"10",x"7f",x"7f",x"13"),
  1876 => (x"67",x"27",x"00",x"00"),
  1877 => (x"39",x"7d",x"45",x"45"),
  1878 => (x"7e",x"3c",x"00",x"00"),
  1879 => (x"30",x"79",x"49",x"4b"),
  1880 => (x"01",x"01",x"00",x"00"),
  1881 => (x"07",x"0f",x"79",x"71"),
  1882 => (x"7f",x"36",x"00",x"00"),
  1883 => (x"36",x"7f",x"49",x"49"),
  1884 => (x"4f",x"06",x"00",x"00"),
  1885 => (x"1e",x"3f",x"69",x"49"),
  1886 => (x"00",x"00",x"00",x"00"),
  1887 => (x"00",x"00",x"66",x"66"),
  1888 => (x"80",x"00",x"00",x"00"),
  1889 => (x"00",x"00",x"66",x"e6"),
  1890 => (x"08",x"08",x"00",x"00"),
  1891 => (x"22",x"22",x"14",x"14"),
  1892 => (x"14",x"14",x"00",x"00"),
  1893 => (x"14",x"14",x"14",x"14"),
  1894 => (x"22",x"22",x"00",x"00"),
  1895 => (x"08",x"08",x"14",x"14"),
  1896 => (x"03",x"02",x"00",x"00"),
  1897 => (x"06",x"0f",x"59",x"51"),
  1898 => (x"41",x"7f",x"3e",x"00"),
  1899 => (x"1e",x"1f",x"55",x"5d"),
  1900 => (x"7f",x"7e",x"00",x"00"),
  1901 => (x"7e",x"7f",x"09",x"09"),
  1902 => (x"7f",x"7f",x"00",x"00"),
  1903 => (x"36",x"7f",x"49",x"49"),
  1904 => (x"3e",x"1c",x"00",x"00"),
  1905 => (x"41",x"41",x"41",x"63"),
  1906 => (x"7f",x"7f",x"00",x"00"),
  1907 => (x"1c",x"3e",x"63",x"41"),
  1908 => (x"7f",x"7f",x"00",x"00"),
  1909 => (x"41",x"41",x"49",x"49"),
  1910 => (x"7f",x"7f",x"00",x"00"),
  1911 => (x"01",x"01",x"09",x"09"),
  1912 => (x"7f",x"3e",x"00",x"00"),
  1913 => (x"7a",x"7b",x"49",x"41"),
  1914 => (x"7f",x"7f",x"00",x"00"),
  1915 => (x"7f",x"7f",x"08",x"08"),
  1916 => (x"41",x"00",x"00",x"00"),
  1917 => (x"00",x"41",x"7f",x"7f"),
  1918 => (x"60",x"20",x"00",x"00"),
  1919 => (x"3f",x"7f",x"40",x"40"),
  1920 => (x"08",x"7f",x"7f",x"00"),
  1921 => (x"41",x"63",x"36",x"1c"),
  1922 => (x"7f",x"7f",x"00",x"00"),
  1923 => (x"40",x"40",x"40",x"40"),
  1924 => (x"06",x"7f",x"7f",x"00"),
  1925 => (x"7f",x"7f",x"06",x"0c"),
  1926 => (x"06",x"7f",x"7f",x"00"),
  1927 => (x"7f",x"7f",x"18",x"0c"),
  1928 => (x"7f",x"3e",x"00",x"00"),
  1929 => (x"3e",x"7f",x"41",x"41"),
  1930 => (x"7f",x"7f",x"00",x"00"),
  1931 => (x"06",x"0f",x"09",x"09"),
  1932 => (x"41",x"7f",x"3e",x"00"),
  1933 => (x"40",x"7e",x"7f",x"61"),
  1934 => (x"7f",x"7f",x"00",x"00"),
  1935 => (x"66",x"7f",x"19",x"09"),
  1936 => (x"6f",x"26",x"00",x"00"),
  1937 => (x"32",x"7b",x"59",x"4d"),
  1938 => (x"01",x"01",x"00",x"00"),
  1939 => (x"01",x"01",x"7f",x"7f"),
  1940 => (x"7f",x"3f",x"00",x"00"),
  1941 => (x"3f",x"7f",x"40",x"40"),
  1942 => (x"3f",x"0f",x"00",x"00"),
  1943 => (x"0f",x"3f",x"70",x"70"),
  1944 => (x"30",x"7f",x"7f",x"00"),
  1945 => (x"7f",x"7f",x"30",x"18"),
  1946 => (x"36",x"63",x"41",x"00"),
  1947 => (x"63",x"36",x"1c",x"1c"),
  1948 => (x"06",x"03",x"01",x"41"),
  1949 => (x"03",x"06",x"7c",x"7c"),
  1950 => (x"59",x"71",x"61",x"01"),
  1951 => (x"41",x"43",x"47",x"4d"),
  1952 => (x"7f",x"00",x"00",x"00"),
  1953 => (x"00",x"41",x"41",x"7f"),
  1954 => (x"06",x"03",x"01",x"00"),
  1955 => (x"60",x"30",x"18",x"0c"),
  1956 => (x"41",x"00",x"00",x"40"),
  1957 => (x"00",x"7f",x"7f",x"41"),
  1958 => (x"06",x"0c",x"08",x"00"),
  1959 => (x"08",x"0c",x"06",x"03"),
  1960 => (x"80",x"80",x"80",x"00"),
  1961 => (x"80",x"80",x"80",x"80"),
  1962 => (x"00",x"00",x"00",x"00"),
  1963 => (x"00",x"04",x"07",x"03"),
  1964 => (x"74",x"20",x"00",x"00"),
  1965 => (x"78",x"7c",x"54",x"54"),
  1966 => (x"7f",x"7f",x"00",x"00"),
  1967 => (x"38",x"7c",x"44",x"44"),
  1968 => (x"7c",x"38",x"00",x"00"),
  1969 => (x"00",x"44",x"44",x"44"),
  1970 => (x"7c",x"38",x"00",x"00"),
  1971 => (x"7f",x"7f",x"44",x"44"),
  1972 => (x"7c",x"38",x"00",x"00"),
  1973 => (x"18",x"5c",x"54",x"54"),
  1974 => (x"7e",x"04",x"00",x"00"),
  1975 => (x"00",x"05",x"05",x"7f"),
  1976 => (x"bc",x"18",x"00",x"00"),
  1977 => (x"7c",x"fc",x"a4",x"a4"),
  1978 => (x"7f",x"7f",x"00",x"00"),
  1979 => (x"78",x"7c",x"04",x"04"),
  1980 => (x"00",x"00",x"00",x"00"),
  1981 => (x"00",x"40",x"7d",x"3d"),
  1982 => (x"80",x"80",x"00",x"00"),
  1983 => (x"00",x"7d",x"fd",x"80"),
  1984 => (x"7f",x"7f",x"00",x"00"),
  1985 => (x"44",x"6c",x"38",x"10"),
  1986 => (x"00",x"00",x"00",x"00"),
  1987 => (x"00",x"40",x"7f",x"3f"),
  1988 => (x"0c",x"7c",x"7c",x"00"),
  1989 => (x"78",x"7c",x"0c",x"18"),
  1990 => (x"7c",x"7c",x"00",x"00"),
  1991 => (x"78",x"7c",x"04",x"04"),
  1992 => (x"7c",x"38",x"00",x"00"),
  1993 => (x"38",x"7c",x"44",x"44"),
  1994 => (x"fc",x"fc",x"00",x"00"),
  1995 => (x"18",x"3c",x"24",x"24"),
  1996 => (x"3c",x"18",x"00",x"00"),
  1997 => (x"fc",x"fc",x"24",x"24"),
  1998 => (x"7c",x"7c",x"00",x"00"),
  1999 => (x"08",x"0c",x"04",x"04"),
  2000 => (x"5c",x"48",x"00",x"00"),
  2001 => (x"20",x"74",x"54",x"54"),
  2002 => (x"3f",x"04",x"00",x"00"),
  2003 => (x"00",x"44",x"44",x"7f"),
  2004 => (x"7c",x"3c",x"00",x"00"),
  2005 => (x"7c",x"7c",x"40",x"40"),
  2006 => (x"3c",x"1c",x"00",x"00"),
  2007 => (x"1c",x"3c",x"60",x"60"),
  2008 => (x"60",x"7c",x"3c",x"00"),
  2009 => (x"3c",x"7c",x"60",x"30"),
  2010 => (x"38",x"6c",x"44",x"00"),
  2011 => (x"44",x"6c",x"38",x"10"),
  2012 => (x"bc",x"1c",x"00",x"00"),
  2013 => (x"1c",x"3c",x"60",x"e0"),
  2014 => (x"64",x"44",x"00",x"00"),
  2015 => (x"44",x"4c",x"5c",x"74"),
  2016 => (x"08",x"08",x"00",x"00"),
  2017 => (x"41",x"41",x"77",x"3e"),
  2018 => (x"00",x"00",x"00",x"00"),
  2019 => (x"00",x"00",x"7f",x"7f"),
  2020 => (x"41",x"41",x"00",x"00"),
  2021 => (x"08",x"08",x"3e",x"77"),
  2022 => (x"01",x"01",x"02",x"00"),
  2023 => (x"01",x"02",x"02",x"03"),
  2024 => (x"7f",x"7f",x"7f",x"00"),
  2025 => (x"7f",x"7f",x"7f",x"7f"),
  2026 => (x"1c",x"08",x"08",x"00"),
  2027 => (x"7f",x"3e",x"3e",x"1c"),
  2028 => (x"3e",x"7f",x"7f",x"7f"),
  2029 => (x"08",x"1c",x"1c",x"3e"),
  2030 => (x"18",x"10",x"00",x"08"),
  2031 => (x"10",x"18",x"7c",x"7c"),
  2032 => (x"30",x"10",x"00",x"00"),
  2033 => (x"10",x"30",x"7c",x"7c"),
  2034 => (x"60",x"30",x"10",x"00"),
  2035 => (x"06",x"1e",x"78",x"60"),
  2036 => (x"3c",x"66",x"42",x"00"),
  2037 => (x"42",x"66",x"3c",x"18"),
  2038 => (x"6a",x"38",x"78",x"00"),
  2039 => (x"38",x"6c",x"c6",x"c2"),
  2040 => (x"00",x"00",x"60",x"00"),
  2041 => (x"60",x"00",x"00",x"60"),
  2042 => (x"5b",x"5e",x"0e",x"00"),
  2043 => (x"1e",x"0e",x"5d",x"5c"),
  2044 => (x"ee",x"c2",x"4c",x"71"),
  2045 => (x"c0",x"4d",x"bf",x"d6"),
  2046 => (x"74",x"1e",x"c0",x"4b"),
  2047 => (x"87",x"c7",x"02",x"ab"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

