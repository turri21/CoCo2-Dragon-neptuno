
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"c0",x"48",x"a6",x"c4"),
     1 => (x"c4",x"87",x"c5",x"78"),
     2 => (x"78",x"c1",x"48",x"a6"),
     3 => (x"73",x"1e",x"66",x"c4"),
     4 => (x"87",x"df",x"ee",x"49"),
     5 => (x"e0",x"c0",x"86",x"c8"),
     6 => (x"87",x"ef",x"ef",x"49"),
     7 => (x"6a",x"4a",x"a5",x"c4"),
     8 => (x"87",x"f0",x"f0",x"49"),
     9 => (x"cb",x"87",x"c6",x"f1"),
    10 => (x"c8",x"83",x"c1",x"85"),
    11 => (x"ff",x"04",x"ab",x"b7"),
    12 => (x"26",x"26",x"87",x"c7"),
    13 => (x"26",x"4c",x"26",x"4d"),
    14 => (x"1e",x"4f",x"26",x"4b"),
    15 => (x"ee",x"c2",x"4a",x"71"),
    16 => (x"ee",x"c2",x"5a",x"da"),
    17 => (x"78",x"c7",x"48",x"da"),
    18 => (x"87",x"dd",x"fe",x"49"),
    19 => (x"73",x"1e",x"4f",x"26"),
    20 => (x"c0",x"4a",x"71",x"1e"),
    21 => (x"d3",x"03",x"aa",x"b7"),
    22 => (x"df",x"ce",x"c2",x"87"),
    23 => (x"87",x"c4",x"05",x"bf"),
    24 => (x"87",x"c2",x"4b",x"c1"),
    25 => (x"ce",x"c2",x"4b",x"c0"),
    26 => (x"87",x"c4",x"5b",x"e3"),
    27 => (x"5a",x"e3",x"ce",x"c2"),
    28 => (x"bf",x"df",x"ce",x"c2"),
    29 => (x"c1",x"9a",x"c1",x"4a"),
    30 => (x"ec",x"49",x"a2",x"c0"),
    31 => (x"48",x"fc",x"87",x"e8"),
    32 => (x"bf",x"df",x"ce",x"c2"),
    33 => (x"87",x"ef",x"fe",x"78"),
    34 => (x"c4",x"4a",x"71",x"1e"),
    35 => (x"49",x"72",x"1e",x"66"),
    36 => (x"26",x"87",x"f5",x"e9"),
    37 => (x"c2",x"1e",x"4f",x"26"),
    38 => (x"49",x"bf",x"df",x"ce"),
    39 => (x"c2",x"87",x"cf",x"e6"),
    40 => (x"e8",x"48",x"ce",x"ee"),
    41 => (x"ee",x"c2",x"78",x"bf"),
    42 => (x"bf",x"ec",x"48",x"ca"),
    43 => (x"ce",x"ee",x"c2",x"78"),
    44 => (x"c3",x"49",x"4a",x"bf"),
    45 => (x"b7",x"c8",x"99",x"ff"),
    46 => (x"71",x"48",x"72",x"2a"),
    47 => (x"d6",x"ee",x"c2",x"b0"),
    48 => (x"0e",x"4f",x"26",x"58"),
    49 => (x"5d",x"5c",x"5b",x"5e"),
    50 => (x"ff",x"4b",x"71",x"0e"),
    51 => (x"ee",x"c2",x"87",x"c8"),
    52 => (x"50",x"c0",x"48",x"c9"),
    53 => (x"f5",x"e5",x"49",x"73"),
    54 => (x"4c",x"49",x"70",x"87"),
    55 => (x"ee",x"cb",x"9c",x"c2"),
    56 => (x"87",x"c3",x"cb",x"49"),
    57 => (x"c2",x"4d",x"49",x"70"),
    58 => (x"bf",x"97",x"c9",x"ee"),
    59 => (x"87",x"e2",x"c1",x"05"),
    60 => (x"c2",x"49",x"66",x"d0"),
    61 => (x"99",x"bf",x"d2",x"ee"),
    62 => (x"d4",x"87",x"d6",x"05"),
    63 => (x"ee",x"c2",x"49",x"66"),
    64 => (x"05",x"99",x"bf",x"ca"),
    65 => (x"49",x"73",x"87",x"cb"),
    66 => (x"70",x"87",x"c3",x"e5"),
    67 => (x"c1",x"c1",x"02",x"98"),
    68 => (x"fe",x"4c",x"c1",x"87"),
    69 => (x"49",x"75",x"87",x"c0"),
    70 => (x"70",x"87",x"d8",x"ca"),
    71 => (x"87",x"c6",x"02",x"98"),
    72 => (x"48",x"c9",x"ee",x"c2"),
    73 => (x"ee",x"c2",x"50",x"c1"),
    74 => (x"05",x"bf",x"97",x"c9"),
    75 => (x"c2",x"87",x"e3",x"c0"),
    76 => (x"49",x"bf",x"d2",x"ee"),
    77 => (x"05",x"99",x"66",x"d0"),
    78 => (x"c2",x"87",x"d6",x"ff"),
    79 => (x"49",x"bf",x"ca",x"ee"),
    80 => (x"05",x"99",x"66",x"d4"),
    81 => (x"73",x"87",x"ca",x"ff"),
    82 => (x"87",x"c2",x"e4",x"49"),
    83 => (x"fe",x"05",x"98",x"70"),
    84 => (x"48",x"74",x"87",x"ff"),
    85 => (x"0e",x"87",x"dc",x"fb"),
    86 => (x"5d",x"5c",x"5b",x"5e"),
    87 => (x"c0",x"86",x"f4",x"0e"),
    88 => (x"bf",x"ec",x"4c",x"4d"),
    89 => (x"48",x"a6",x"c4",x"7e"),
    90 => (x"bf",x"d6",x"ee",x"c2"),
    91 => (x"c0",x"1e",x"c1",x"78"),
    92 => (x"fd",x"49",x"c7",x"1e"),
    93 => (x"86",x"c8",x"87",x"cd"),
    94 => (x"cd",x"02",x"98",x"70"),
    95 => (x"fb",x"49",x"ff",x"87"),
    96 => (x"da",x"c1",x"87",x"cc"),
    97 => (x"87",x"c6",x"e3",x"49"),
    98 => (x"ee",x"c2",x"4d",x"c1"),
    99 => (x"02",x"bf",x"97",x"c9"),
   100 => (x"fe",x"d4",x"87",x"c3"),
   101 => (x"ce",x"ee",x"c2",x"87"),
   102 => (x"ce",x"c2",x"4b",x"bf"),
   103 => (x"c0",x"05",x"bf",x"df"),
   104 => (x"fd",x"c3",x"87",x"e9"),
   105 => (x"87",x"e6",x"e2",x"49"),
   106 => (x"e2",x"49",x"fa",x"c3"),
   107 => (x"49",x"73",x"87",x"e0"),
   108 => (x"71",x"99",x"ff",x"c3"),
   109 => (x"fb",x"49",x"c0",x"1e"),
   110 => (x"49",x"73",x"87",x"ce"),
   111 => (x"71",x"29",x"b7",x"c8"),
   112 => (x"fb",x"49",x"c1",x"1e"),
   113 => (x"86",x"c8",x"87",x"c2"),
   114 => (x"c2",x"87",x"fa",x"c5"),
   115 => (x"4b",x"bf",x"d2",x"ee"),
   116 => (x"87",x"dd",x"02",x"9b"),
   117 => (x"bf",x"db",x"ce",x"c2"),
   118 => (x"87",x"d7",x"c7",x"49"),
   119 => (x"c4",x"05",x"98",x"70"),
   120 => (x"d2",x"4b",x"c0",x"87"),
   121 => (x"49",x"e0",x"c2",x"87"),
   122 => (x"c2",x"87",x"fc",x"c6"),
   123 => (x"c6",x"58",x"df",x"ce"),
   124 => (x"db",x"ce",x"c2",x"87"),
   125 => (x"73",x"78",x"c0",x"48"),
   126 => (x"05",x"99",x"c2",x"49"),
   127 => (x"eb",x"c3",x"87",x"cd"),
   128 => (x"87",x"ca",x"e1",x"49"),
   129 => (x"99",x"c2",x"49",x"70"),
   130 => (x"fb",x"87",x"c2",x"02"),
   131 => (x"c1",x"49",x"73",x"4c"),
   132 => (x"87",x"cd",x"05",x"99"),
   133 => (x"e0",x"49",x"f4",x"c3"),
   134 => (x"49",x"70",x"87",x"f4"),
   135 => (x"c2",x"02",x"99",x"c2"),
   136 => (x"73",x"4c",x"fa",x"87"),
   137 => (x"05",x"99",x"c8",x"49"),
   138 => (x"f5",x"c3",x"87",x"cd"),
   139 => (x"87",x"de",x"e0",x"49"),
   140 => (x"99",x"c2",x"49",x"70"),
   141 => (x"c2",x"87",x"d4",x"02"),
   142 => (x"02",x"bf",x"da",x"ee"),
   143 => (x"c1",x"48",x"87",x"c9"),
   144 => (x"de",x"ee",x"c2",x"88"),
   145 => (x"ff",x"87",x"c2",x"58"),
   146 => (x"73",x"4d",x"c1",x"4c"),
   147 => (x"05",x"99",x"c4",x"49"),
   148 => (x"f2",x"c3",x"87",x"ce"),
   149 => (x"f5",x"df",x"ff",x"49"),
   150 => (x"c2",x"49",x"70",x"87"),
   151 => (x"87",x"db",x"02",x"99"),
   152 => (x"bf",x"da",x"ee",x"c2"),
   153 => (x"b7",x"c7",x"48",x"7e"),
   154 => (x"87",x"cb",x"03",x"a8"),
   155 => (x"80",x"c1",x"48",x"6e"),
   156 => (x"58",x"de",x"ee",x"c2"),
   157 => (x"fe",x"87",x"c2",x"c0"),
   158 => (x"c3",x"4d",x"c1",x"4c"),
   159 => (x"df",x"ff",x"49",x"fd"),
   160 => (x"49",x"70",x"87",x"cc"),
   161 => (x"d5",x"02",x"99",x"c2"),
   162 => (x"da",x"ee",x"c2",x"87"),
   163 => (x"c9",x"c0",x"02",x"bf"),
   164 => (x"da",x"ee",x"c2",x"87"),
   165 => (x"c0",x"78",x"c0",x"48"),
   166 => (x"4c",x"fd",x"87",x"c2"),
   167 => (x"fa",x"c3",x"4d",x"c1"),
   168 => (x"e9",x"de",x"ff",x"49"),
   169 => (x"c2",x"49",x"70",x"87"),
   170 => (x"87",x"d9",x"02",x"99"),
   171 => (x"bf",x"da",x"ee",x"c2"),
   172 => (x"a8",x"b7",x"c7",x"48"),
   173 => (x"87",x"c9",x"c0",x"03"),
   174 => (x"48",x"da",x"ee",x"c2"),
   175 => (x"c2",x"c0",x"78",x"c7"),
   176 => (x"c1",x"4c",x"fc",x"87"),
   177 => (x"ac",x"b7",x"c0",x"4d"),
   178 => (x"87",x"d1",x"c0",x"03"),
   179 => (x"c1",x"4a",x"66",x"c4"),
   180 => (x"02",x"6a",x"82",x"d8"),
   181 => (x"6a",x"87",x"c6",x"c0"),
   182 => (x"73",x"49",x"74",x"4b"),
   183 => (x"c3",x"1e",x"c0",x"0f"),
   184 => (x"da",x"c1",x"1e",x"f0"),
   185 => (x"87",x"db",x"f7",x"49"),
   186 => (x"98",x"70",x"86",x"c8"),
   187 => (x"87",x"e2",x"c0",x"02"),
   188 => (x"c2",x"48",x"a6",x"c8"),
   189 => (x"78",x"bf",x"da",x"ee"),
   190 => (x"cb",x"49",x"66",x"c8"),
   191 => (x"48",x"66",x"c4",x"91"),
   192 => (x"7e",x"70",x"80",x"71"),
   193 => (x"c0",x"02",x"bf",x"6e"),
   194 => (x"bf",x"6e",x"87",x"c8"),
   195 => (x"49",x"66",x"c8",x"4b"),
   196 => (x"9d",x"75",x"0f",x"73"),
   197 => (x"87",x"c8",x"c0",x"02"),
   198 => (x"bf",x"da",x"ee",x"c2"),
   199 => (x"87",x"c9",x"f3",x"49"),
   200 => (x"bf",x"e3",x"ce",x"c2"),
   201 => (x"87",x"dd",x"c0",x"02"),
   202 => (x"87",x"c7",x"c2",x"49"),
   203 => (x"c0",x"02",x"98",x"70"),
   204 => (x"ee",x"c2",x"87",x"d3"),
   205 => (x"f2",x"49",x"bf",x"da"),
   206 => (x"49",x"c0",x"87",x"ef"),
   207 => (x"c2",x"87",x"cf",x"f4"),
   208 => (x"c0",x"48",x"e3",x"ce"),
   209 => (x"f3",x"8e",x"f4",x"78"),
   210 => (x"5e",x"0e",x"87",x"e9"),
   211 => (x"0e",x"5d",x"5c",x"5b"),
   212 => (x"c2",x"4c",x"71",x"1e"),
   213 => (x"49",x"bf",x"d6",x"ee"),
   214 => (x"4d",x"a1",x"cd",x"c1"),
   215 => (x"69",x"81",x"d1",x"c1"),
   216 => (x"02",x"9c",x"74",x"7e"),
   217 => (x"a5",x"c4",x"87",x"cf"),
   218 => (x"c2",x"7b",x"74",x"4b"),
   219 => (x"49",x"bf",x"d6",x"ee"),
   220 => (x"6e",x"87",x"c8",x"f3"),
   221 => (x"05",x"9c",x"74",x"7b"),
   222 => (x"4b",x"c0",x"87",x"c4"),
   223 => (x"4b",x"c1",x"87",x"c2"),
   224 => (x"c9",x"f3",x"49",x"73"),
   225 => (x"02",x"66",x"d4",x"87"),
   226 => (x"da",x"49",x"87",x"c7"),
   227 => (x"c2",x"4a",x"70",x"87"),
   228 => (x"c2",x"4a",x"c0",x"87"),
   229 => (x"26",x"5a",x"e7",x"ce"),
   230 => (x"00",x"87",x"d8",x"f2"),
   231 => (x"00",x"00",x"00",x"00"),
   232 => (x"00",x"00",x"00",x"00"),
   233 => (x"1e",x"00",x"00",x"00"),
   234 => (x"c8",x"ff",x"4a",x"71"),
   235 => (x"a1",x"72",x"49",x"bf"),
   236 => (x"1e",x"4f",x"26",x"48"),
   237 => (x"89",x"bf",x"c8",x"ff"),
   238 => (x"c0",x"c0",x"c0",x"fe"),
   239 => (x"01",x"a9",x"c0",x"c0"),
   240 => (x"4a",x"c0",x"87",x"c4"),
   241 => (x"4a",x"c1",x"87",x"c2"),
   242 => (x"4f",x"26",x"48",x"72"),
   243 => (x"5c",x"5b",x"5e",x"0e"),
   244 => (x"4b",x"71",x"0e",x"5d"),
   245 => (x"d0",x"4c",x"d4",x"ff"),
   246 => (x"78",x"c0",x"48",x"66"),
   247 => (x"db",x"ff",x"49",x"d6"),
   248 => (x"ff",x"c3",x"87",x"ec"),
   249 => (x"c3",x"49",x"6c",x"7c"),
   250 => (x"4d",x"71",x"99",x"ff"),
   251 => (x"99",x"f0",x"c3",x"49"),
   252 => (x"05",x"a9",x"e0",x"c1"),
   253 => (x"ff",x"c3",x"87",x"cb"),
   254 => (x"c3",x"48",x"6c",x"7c"),
   255 => (x"08",x"66",x"d0",x"98"),
   256 => (x"7c",x"ff",x"c3",x"78"),
   257 => (x"c8",x"49",x"4a",x"6c"),
   258 => (x"7c",x"ff",x"c3",x"31"),
   259 => (x"b2",x"71",x"4a",x"6c"),
   260 => (x"31",x"c8",x"49",x"72"),
   261 => (x"6c",x"7c",x"ff",x"c3"),
   262 => (x"72",x"b2",x"71",x"4a"),
   263 => (x"c3",x"31",x"c8",x"49"),
   264 => (x"4a",x"6c",x"7c",x"ff"),
   265 => (x"d0",x"ff",x"b2",x"71"),
   266 => (x"78",x"e0",x"c0",x"48"),
   267 => (x"c2",x"02",x"9b",x"73"),
   268 => (x"75",x"7b",x"72",x"87"),
   269 => (x"26",x"4d",x"26",x"48"),
   270 => (x"26",x"4b",x"26",x"4c"),
   271 => (x"4f",x"26",x"1e",x"4f"),
   272 => (x"5c",x"5b",x"5e",x"0e"),
   273 => (x"76",x"86",x"f8",x"0e"),
   274 => (x"49",x"a6",x"c8",x"1e"),
   275 => (x"c4",x"87",x"fd",x"fd"),
   276 => (x"6e",x"4b",x"70",x"86"),
   277 => (x"03",x"a8",x"c2",x"48"),
   278 => (x"73",x"87",x"c6",x"c3"),
   279 => (x"9a",x"f0",x"c3",x"4a"),
   280 => (x"02",x"aa",x"d0",x"c1"),
   281 => (x"e0",x"c1",x"87",x"c7"),
   282 => (x"f4",x"c2",x"05",x"aa"),
   283 => (x"c8",x"49",x"73",x"87"),
   284 => (x"87",x"c3",x"02",x"99"),
   285 => (x"73",x"87",x"c6",x"ff"),
   286 => (x"c2",x"9c",x"c3",x"4c"),
   287 => (x"cd",x"c1",x"05",x"ac"),
   288 => (x"49",x"66",x"c4",x"87"),
   289 => (x"1e",x"71",x"31",x"c9"),
   290 => (x"d4",x"4a",x"66",x"c4"),
   291 => (x"de",x"ee",x"c2",x"92"),
   292 => (x"fe",x"81",x"72",x"49"),
   293 => (x"c4",x"87",x"d8",x"d4"),
   294 => (x"c0",x"1e",x"49",x"66"),
   295 => (x"d9",x"ff",x"49",x"e3"),
   296 => (x"49",x"d8",x"87",x"d1"),
   297 => (x"87",x"e6",x"d8",x"ff"),
   298 => (x"c2",x"1e",x"c0",x"c8"),
   299 => (x"fd",x"49",x"ce",x"dd"),
   300 => (x"ff",x"87",x"e8",x"f0"),
   301 => (x"e0",x"c0",x"48",x"d0"),
   302 => (x"ce",x"dd",x"c2",x"78"),
   303 => (x"4a",x"66",x"d0",x"1e"),
   304 => (x"ee",x"c2",x"92",x"d4"),
   305 => (x"81",x"72",x"49",x"de"),
   306 => (x"87",x"e0",x"d2",x"fe"),
   307 => (x"ac",x"c1",x"86",x"d0"),
   308 => (x"87",x"cd",x"c1",x"05"),
   309 => (x"c9",x"49",x"66",x"c4"),
   310 => (x"c4",x"1e",x"71",x"31"),
   311 => (x"92",x"d4",x"4a",x"66"),
   312 => (x"49",x"de",x"ee",x"c2"),
   313 => (x"d3",x"fe",x"81",x"72"),
   314 => (x"dd",x"c2",x"87",x"c5"),
   315 => (x"66",x"c8",x"1e",x"ce"),
   316 => (x"c2",x"92",x"d4",x"4a"),
   317 => (x"72",x"49",x"de",x"ee"),
   318 => (x"ec",x"d0",x"fe",x"81"),
   319 => (x"49",x"66",x"c8",x"87"),
   320 => (x"49",x"e3",x"c0",x"1e"),
   321 => (x"87",x"eb",x"d7",x"ff"),
   322 => (x"d7",x"ff",x"49",x"d7"),
   323 => (x"c0",x"c8",x"87",x"c0"),
   324 => (x"ce",x"dd",x"c2",x"1e"),
   325 => (x"ec",x"ee",x"fd",x"49"),
   326 => (x"ff",x"86",x"d0",x"87"),
   327 => (x"e0",x"c0",x"48",x"d0"),
   328 => (x"fc",x"8e",x"f8",x"78"),
   329 => (x"5e",x"0e",x"87",x"d1"),
   330 => (x"0e",x"5d",x"5c",x"5b"),
   331 => (x"ff",x"4d",x"71",x"1e"),
   332 => (x"66",x"d4",x"4c",x"d4"),
   333 => (x"b7",x"c3",x"48",x"7e"),
   334 => (x"87",x"c5",x"06",x"a8"),
   335 => (x"e2",x"c1",x"48",x"c0"),
   336 => (x"fe",x"49",x"75",x"87"),
   337 => (x"75",x"87",x"f9",x"e0"),
   338 => (x"4b",x"66",x"c4",x"1e"),
   339 => (x"ee",x"c2",x"93",x"d4"),
   340 => (x"49",x"73",x"83",x"de"),
   341 => (x"87",x"f5",x"cb",x"fe"),
   342 => (x"4b",x"6b",x"83",x"c8"),
   343 => (x"c8",x"48",x"d0",x"ff"),
   344 => (x"7c",x"dd",x"78",x"e1"),
   345 => (x"ff",x"c3",x"49",x"73"),
   346 => (x"73",x"7c",x"71",x"99"),
   347 => (x"29",x"b7",x"c8",x"49"),
   348 => (x"71",x"99",x"ff",x"c3"),
   349 => (x"d0",x"49",x"73",x"7c"),
   350 => (x"ff",x"c3",x"29",x"b7"),
   351 => (x"73",x"7c",x"71",x"99"),
   352 => (x"29",x"b7",x"d8",x"49"),
   353 => (x"7c",x"c0",x"7c",x"71"),
   354 => (x"7c",x"7c",x"7c",x"7c"),
   355 => (x"7c",x"7c",x"7c",x"7c"),
   356 => (x"c0",x"7c",x"7c",x"7c"),
   357 => (x"66",x"c4",x"78",x"e0"),
   358 => (x"ff",x"49",x"dc",x"1e"),
   359 => (x"c8",x"87",x"d4",x"d5"),
   360 => (x"26",x"48",x"73",x"86"),
   361 => (x"0e",x"87",x"ce",x"fa"),
   362 => (x"5d",x"5c",x"5b",x"5e"),
   363 => (x"7e",x"71",x"1e",x"0e"),
   364 => (x"6e",x"4b",x"d4",x"ff"),
   365 => (x"c6",x"ef",x"c2",x"1e"),
   366 => (x"d0",x"ca",x"fe",x"49"),
   367 => (x"70",x"86",x"c4",x"87"),
   368 => (x"c3",x"02",x"9d",x"4d"),
   369 => (x"ef",x"c2",x"87",x"c3"),
   370 => (x"6e",x"4c",x"bf",x"ce"),
   371 => (x"ef",x"de",x"fe",x"49"),
   372 => (x"48",x"d0",x"ff",x"87"),
   373 => (x"c1",x"78",x"c5",x"c8"),
   374 => (x"4a",x"c0",x"7b",x"d6"),
   375 => (x"82",x"c1",x"7b",x"15"),
   376 => (x"aa",x"b7",x"e0",x"c0"),
   377 => (x"ff",x"87",x"f5",x"04"),
   378 => (x"78",x"c4",x"48",x"d0"),
   379 => (x"c1",x"78",x"c5",x"c8"),
   380 => (x"7b",x"c1",x"7b",x"d3"),
   381 => (x"9c",x"74",x"78",x"c4"),
   382 => (x"87",x"fc",x"c1",x"02"),
   383 => (x"7e",x"ce",x"dd",x"c2"),
   384 => (x"8c",x"4d",x"c0",x"c8"),
   385 => (x"03",x"ac",x"b7",x"c0"),
   386 => (x"c0",x"c8",x"87",x"c6"),
   387 => (x"4c",x"c0",x"4d",x"a4"),
   388 => (x"97",x"ff",x"e9",x"c2"),
   389 => (x"99",x"d0",x"49",x"bf"),
   390 => (x"c0",x"87",x"d2",x"02"),
   391 => (x"c6",x"ef",x"c2",x"1e"),
   392 => (x"c4",x"cc",x"fe",x"49"),
   393 => (x"70",x"86",x"c4",x"87"),
   394 => (x"ef",x"c0",x"4a",x"49"),
   395 => (x"ce",x"dd",x"c2",x"87"),
   396 => (x"c6",x"ef",x"c2",x"1e"),
   397 => (x"f0",x"cb",x"fe",x"49"),
   398 => (x"70",x"86",x"c4",x"87"),
   399 => (x"d0",x"ff",x"4a",x"49"),
   400 => (x"78",x"c5",x"c8",x"48"),
   401 => (x"6e",x"7b",x"d4",x"c1"),
   402 => (x"6e",x"7b",x"bf",x"97"),
   403 => (x"70",x"80",x"c1",x"48"),
   404 => (x"05",x"8d",x"c1",x"7e"),
   405 => (x"ff",x"87",x"f0",x"ff"),
   406 => (x"78",x"c4",x"48",x"d0"),
   407 => (x"c5",x"05",x"9a",x"72"),
   408 => (x"c0",x"48",x"c0",x"87"),
   409 => (x"1e",x"c1",x"87",x"e5"),
   410 => (x"49",x"c6",x"ef",x"c2"),
   411 => (x"87",x"d8",x"c9",x"fe"),
   412 => (x"9c",x"74",x"86",x"c4"),
   413 => (x"87",x"c4",x"fe",x"05"),
   414 => (x"c8",x"48",x"d0",x"ff"),
   415 => (x"d3",x"c1",x"78",x"c5"),
   416 => (x"c4",x"7b",x"c0",x"7b"),
   417 => (x"c2",x"48",x"c1",x"78"),
   418 => (x"26",x"48",x"c0",x"87"),
   419 => (x"4c",x"26",x"4d",x"26"),
   420 => (x"4f",x"26",x"4b",x"26"),
   421 => (x"5c",x"5b",x"5e",x"0e"),
   422 => (x"cc",x"4b",x"71",x"0e"),
   423 => (x"87",x"d8",x"02",x"66"),
   424 => (x"8c",x"f0",x"c0",x"4c"),
   425 => (x"74",x"87",x"d8",x"02"),
   426 => (x"02",x"8a",x"c1",x"4a"),
   427 => (x"02",x"8a",x"87",x"d1"),
   428 => (x"02",x"8a",x"87",x"cd"),
   429 => (x"87",x"d7",x"87",x"c9"),
   430 => (x"ea",x"fb",x"49",x"73"),
   431 => (x"74",x"87",x"d0",x"87"),
   432 => (x"f9",x"49",x"c0",x"1e"),
   433 => (x"1e",x"74",x"87",x"e0"),
   434 => (x"d9",x"f9",x"49",x"73"),
   435 => (x"fe",x"86",x"c8",x"87"),
   436 => (x"1e",x"00",x"87",x"fc"),
   437 => (x"bf",x"e1",x"dc",x"c2"),
   438 => (x"c2",x"b9",x"c1",x"49"),
   439 => (x"ff",x"59",x"e5",x"dc"),
   440 => (x"ff",x"c3",x"48",x"d4"),
   441 => (x"48",x"d0",x"ff",x"78"),
   442 => (x"ff",x"78",x"e1",x"c8"),
   443 => (x"78",x"c1",x"48",x"d4"),
   444 => (x"78",x"71",x"31",x"c4"),
   445 => (x"c0",x"48",x"d0",x"ff"),
   446 => (x"4f",x"26",x"78",x"e0"),
   447 => (x"d5",x"dc",x"c2",x"1e"),
   448 => (x"c6",x"ef",x"c2",x"1e"),
   449 => (x"c4",x"c5",x"fe",x"49"),
   450 => (x"70",x"86",x"c4",x"87"),
   451 => (x"87",x"c3",x"02",x"98"),
   452 => (x"26",x"87",x"c0",x"ff"),
   453 => (x"4b",x"35",x"31",x"4f"),
   454 => (x"20",x"20",x"5a",x"48"),
   455 => (x"47",x"46",x"43",x"20"),
   456 => (x"00",x"00",x"00",x"00"),
   457 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

